XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����`�rd��߇R�(W����y��Ňw`���g�L$��;'���(!0�P�M���4�&]�w荏����%fG:��
�;�����+ _���wa�X�3T�c�Dr�����y&��(p��80u�(�83�EK�� �;� ��

��v�۸vT����$>�Q;�mTvjݘ*KJ���|ޗ�V�?p���K�3\ť����]��gm��S߱A�>5�K�92 RF����t�k�`RirL$���vz���e>̧Fc �,l�r�c˜�*�x
�w��:yGai�� I,�UK,��ߖ�[\ǫU�=�����o�Hy
r����R�|Q%������!fhY��>V}p��[)���|�ʩ���%�$GfbY����`�軃�����3�_1�����V�f���t�(���iSe_f�Dn3��YxԵ.#���כ��F�[���bѠ��i��-E@�.�c4��ٶK�{��E\u/q�lnE�w��-i����[��H۹m�h������ެ7!�ի���_�7���b.�k��\���S�V]O�?��s"m�1����K��h4&�/tۘj�5z���NT#[iӮJ�]e=��i*�ˋ�'����U��?&���`mx}ާ�C����'�l���i\�w��9�HB�ޘ�R�A�n|��D���s��M�<y�qs<A���!�|
l�|&�W�AA!Ҥ=��ZO7�)�x����Gs�����r):���9ᄊ��p,�XlxVHYEB    1602     7a0��]���I�T���]���91�P~����$��mA��/"���)��(��bH|/M����O����Rp�5��b]��e��Z54�<F�	-r���o4�T��YZ�s������#%��Pz��[�~ק��pO~��Y�Dh#�w��	箴k��@Xc�@wL�Բ��tK��?����?w�D���pS�[.�ǝ����g�������K~�f�"��N9.XĻÂ�fF{z���I�L�y�po���^J�6����W�@����$ت!.��v߆����v�E@>�q����4���J4W'q�O:����TH����<x��A�"�[��xs�so��Vjw��7_�p�C)����$:�%l'��Z��P����'җ=� �:��;��^�S���(�K��]�7<a�ls�KS�@�HJ�u�	�	�`L�E�����x>�AM�ź�M�5�
�B$Z`U�f_P�rU���\S��3�Ң4��n��\��ϋN�� ��#���͜u*P��NVSG���������Z\۪�X(2��#v���/iU^M0�/�%z��5��D��[p5u.�3���e���>`J����Nx"��4[�b��w��%f`w0��F��z=h��lJ}K#�)D��2.���I�bKxO���~S�$�Q�nAx��}=����C��s����T�e)(s���dM���N�ׯ�9��y^Oh �;�ݴ3XOOQ�Y�e;�~#���	L�r��Y
 �䁱���9�И:Jé����K;t<_�q�`_��/奩I����!��;�f�]��/�(e��|$����i�9�������=zo{k;1�!Q�]MΤ�L?���'�2&y�E`���	�0������^i+-E�D�\j�j��m����Q@e���ƀ�C%ϻ�앶J�Xо���w���a7i�qk��q�_#�-�`^㈐�t͞,x�孲9$;�{�@��gfw���両Cϋu���a��c�e�`�C���)x��ւݦ�WU{{�&�+&��_x&��_M��O#k.cYp���[��F :�dP_	Q@��hj7�i�Z�Y��Ю� R����߁UѴ6�>�=Lu���I�^�����k��ƕC�&����[��T���V��k�{IsUp�K��@N< =^R��;��P�U+1�Q�'��6���C.*)y�=��S	��ެ���}�m���u���(u"U"Y���*���4/���- ����y��%��	����j�� �v��x�KE���{5��M>��O~�s��Ɯ�<~s�� �A�r<8����C(��+r����4ڴ�mF�2��]�n���܆��	�؝#�L�(W) d�r�ᚿ��^96��މ������8�*X:�l����dö$�MʍF��H܊ �u�K�W����i�R�Y�)q�xԖ������oK�V�P�Eěj�,p��b[��n�X7N��%��ZL�k|��a��0�����L�
$^�
�j5��U��ɠ;ZV�Dy%���+<Y�_iQ����b�����=�AUwE}�+hɰ4�9�J8�[9�F�yٵ0��0Ѻ3�j,J\�s~n���u��/ʌ�Z����;E`�Tr�� ��KؕjQ�����U�ZBG�!�_� {�`�4vG��N����� d[����q-P����T�F]M[v�d׽�c��Yi�j
]�I���ƨI�%��#ꛝ$����u;���J]�B�Wo���q��Q�vt�g�&9��WkA���	�"D�U������LFQ��r���͔�pXG߾������J]a��cgV�=_�8�0�c�^]y�r��CNJ�`��g�ƌ�f�J���J#Y������|���jA��(�I�fi���ME4L����H2�ڿ�`j�*�l:�A��m�Xׄ��߻;��+�2�6