XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Y�2��6^�I].�b(2�K���H�խ���̨������xܲ��:�3��s�4 �y�ֶ]����L�Z��D�̲mCҮ�c��WЀ\���E�Θ5��w�������)ޤ������
G��1��]Z�1����Ou^�>a��J��{��岛Tm�q�o"����Q�W�?4 N�P����_�[���Ov@�j��2Wj������^��N�u
�It��<K����i��ZN ������rLQ�Rv���`���o��:I�2.��hJL"1��č<F �ajÈ�9%xEh������ R�b4q.6�#��Ħ7F�����vmHs���Wϡ�f���C�5���;�_��pr�&�d�c�e����$J�65U�3���*�(|���±&i���%��z@/��ߎ5F5X��n��]~8��5�f����2eð�YTV,Ϸ��S�UA�s�B���HizT�3�Lν`f��.U�n�H+���R�0��'/G��
�����6�\<b����ڟ�����2	�gN�`�$�;\BH���|gm��Y��������7�	��s�K�"�gBD��U~vF->j�#��e
��*@jooڛ��N8�ֺ�c%��}'���D���D	�}֨&�Ŗ"��U�����S�v6�X���)q=Ŭ��n�xp0ɒ���o��E�m�b4P,���*�P��3��E��2���녽�ֲO�F��((w#|�A��Şy!G� �Z����V{%�+(�XlxVHYEB    3189     890~�bg�,m����X~�ͻ��{=��S2�e��`fLOGӅ }�Ë�t���K��_40*a�W�Y������P���?f�v�Q�����i��d��X�ε�2�Kk-�t�$w�36Ay`��-�#Oc(Y	�&��=�P7ֳrh��sn| ���}+�\��Y�?����Sv�K���{xzQ�#��.��#C� ܤ� �̂��71�P\7#B����?#C�۷� _ۉ���-�Rh�1g&_���؜���-?�e�Ð��u,BV�������T��1�Ϛ��7�2q \�t��IR�b[5q�ȿ�3o}�s�ڬ��v�˩3�����N��3�a�x#�����R�^9�|���m^�͹݊�E�t͕E�~D��/�)�\�dU����IJ�5�:�v�*���M�d��3رT��V���D�CD�3 ѳ�P@ָ�al�+Ԓ���8��O����a��B��V.��p��,��&kpKg�����T�̣
��|V[�����E|i�f4;���w��+�����įXx��R5���\��I�5��v��yV�J??�de&�j빪�-�t'���ة}7J�q�,u�*�u�vQ�ە�'9p����,��QS� ����53�ň`Հ���j�� YzI��9�t�ҦC�zh��N�$q]���39��4�Ƙ�Lz��̾�1���*뇈����}�'�9��O@/)����]�du����}͌8���3� �W���!J��\��J���;�G�x�K���"��^�����N�k���`��t�Ɵt)Z��n��X+�"�}�|��֣�`X�����W��a���W������uN�����M-��!V�8�&64^��+XN29�%�W�O%��@�Y�JAghQ��|� �&�כ�~z-@w�����lo�Z�[�5����G!	*��:�#���P�B�nQN��K��"��s/'��򙦜Y���&�����(��V�. BF nJ5�3Gd��3Z�TY(���>�M/v�\�xH\t]�_Mx��dq�Q�;!!��꾹QѠC.ɭ��O-$�&�w���LR�q�l�[u�	Pb�>�!b�$�A0v	P^N��NoC+�(��F����� �ی�c�a�#���ZTC���N4Z�` ҢA�&��$����C%c6��Êr��`(p��Hl�لsvz��펊o�s�_�Ķ(��yA�$��P[�{yʢ�R:xf?������qd{a�46�|�e��N���y���^@ݲ�COU��yB����hc`!N��"T_����'-��"c4[�xNc� L%2���W.�r�Ÿ�fp-s�����,�)-c��80dfK3���:�|���χbb�m�lbZ�~IGV��t�4Ț�_`�kb)��w���ߪ��Mr�8o���/�ȣT���fL��2z��j$_e&�%PCc*�_�:�`� \s�/}���.L6�5"�Bmc��� ��*��\᰾!!��J+�dϷt��)򛭻�L�N)���l�p�t��͖�̣�٩˖��Oħ��&v�N"cD�0N�� ��u76ox,��s���~������8���2~�h�l�E�O�d͈�^��ެ����F/�,����e`4Tlt�����GS�$��?�!�������Ƙwu�$M��?����V���7c+$�K�z�����fs7%�H$�h>�Q����Fڰ�O�������7r��%���C��yy_
N7�:;`�X��XB��ԝ|?�M��S�K�|=�� s�.�������.?W�^���}��(l+$�D���Q��s�J�����?/�K;����=I�@}���>ŐXk-F�\J����@�[�����0�y����N�?�n
��Pז��z��q&��}�A'[�����.�����3`RwBPi�w(��&����������4ů2�>����r��� Q���=z�pQaq�\��BL�jS_��.�Hk�ߞ��0lA�^��3sKV�c��̵�i�
wL���1���U%ֹ6AT�\����Ťק ��l�z~�4��\_1wm�ɳa�)ѰnO#7����`�e���>�W&�kA�]̀����}$�BN]�v� ]��z����*i3��T�ѷ
��S�.80��q��*��v��>���sM�����+�]�Ȥ\���.�