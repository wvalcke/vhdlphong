XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ta�(FSك{�bM�S�
b�ƙ�"WX�l��5`�uČ1�0���d�T��u�y�_��߀�l���t!'��uEܹRRu����c�oi[���.J�uz?F�~���u����	��U}��Ç��'{���H$���h�m�K_!M54���t��ШO��h���'0f����l�P��^s(�YMaj��W��`px»%tޱg=�]�j� $���J�i8��� �J�������+�D�\���g�`-��vfq��|�0�MŅ�#�%Z��͏�T���a�&�yۈ��;�;��`OmQb$`�s�9r�?x��5T��J���;���i��=HO�����8�������U_�mF�L�	�&�-��0�E�+a�ySSM����P���f�:Og���9�\-nuz�h3���![,X�����-��nгw�����H'C��J*z��L��!�L���ʿ�>�YmdN�~��_p��Հ���]��8�B{7;5��2E�t��V�GcLk�)j��w��14d^��/6��ɸ�yo.Okfo�`�_�%�z9a�e�ܫ��56-�*K�zu��^'Tw׷'���P�&:pcը�$ϐH�a�ҵqŐ��gʤv��:�y��2�-��Z༌�R����N���t�~���ɓ�2��e�c�(اt�B�$�?R�V|/��:���`Cn(ӭ�R6����dQs>i�͉��p"�>}F���;1�W�1m ʶ��G���E���E����OP�$Z�r)�ga�����p�6ǾF>��XlxVHYEB    5ee8    14d0��B4~��a�,�Qa'#kA#?�1��
Fiq�����Zh�diiz*峬�͔7�=�Y��@���v/�CWr��
�iDqv��&�dW(���Opm�]��H\1�H_���j�W4���:�s����0Uěc�����d.��.C6��{̭��_E���K��H��L̑W�]u�[5���&�sWp�k>3�v���|�Cv��H�@�h����]��Ǆ|���,���ker���ڂj鬾�������O�tu����];0c���{�^k�qE��`�����o3�X��S	�4��:,���`@;���Я"-���Ϧ��_"�0��ի�a���I���J11'#b#z�;�M��(bjiV�c�����]��KL��o��.y�N��>��i�<K~���,���n���� g�D-��$������
��Ϋy�q�9�lwvX�/�Md�6��⭥�v��a%���1��K�T�f�}����xv�.RB��O;E[σ�+0�**M,2e�L��<���m3d������S�W�'��v_��|ϲ�\v	i ���b��ێ���[B��J�������]��Z��>��sR1�y�|�(1�B�"/��,Ϟ�_|�]�~1#��MO��߰�ys�����`H�eeI�ȁʖ��t����w;G�a#�^���L�����O�vh�A�-��������9��hc7/�����PL����S� $����Q��9j��E�+����N6�*���6�m��f��ӣI��[�/7��q4w�R�mv�>�ꋃ-�1�к�Ծݙ;�,���b�����Zq�"{{���Y%��|
DU3�K�V0�|�,�|%q�& ���V`�|�+B��g�=�ҡot��b��ֈ�[
��<�Z%����>x��M����声sobCo�翶>��-�	�ݎ� `cՑ�kﭴ��7S�؃Z�W�ف�`>�)�2���W�8"-�B5��bJ�Y���E���_q���,��R��L1���n����>�
v�%H���i�es�5��
���;����zL�)(�7U�|���:�T�mby��o<<ɀ��2�"�#�m,��=�R��;j!������C`��Yy�~����b������|��9Ykx��u�� �<C�X5������|����0���&���e�DLؐ��U��K"��,�IEy�ޭv�2@��6�4�4�45RsiV�l��~_Ǆ��@�984�b�z9C
�!m,KＮͅbl��	O=�Qx�o,W�C�4Z;G��^��\KSb�Z��M
:�Z�"*�4xT:f�[;�hڪ.(o�S��[!m,qQ*j��|����>��C_m���iq�\�~���@sta��\T������ͺ|���t<_4���oF��Ϝc3�sM�1�ݲ�AX�ƅ-V�[׹�( $���RNXE:Jg����d�ۓ@ia�q�}[ 
SG�����x����
��S�iߢ Aß����G����.%rD��o��p�<�d�]��C�q���y��$tPss%�nU�2�㾷 '�tˊ�K�j��hM��q�*�m���x�q����/���b^45PI���.?����O|�3����c�e���P�����i�U��1G��}���(1vODmG�*Bsɫ��"�$E5)��kI������F���Z�yI3��ĩ|�D�q�\c�Z�q{#���7��M�
��a9�\�TR�NZ��X��l����u�SH�#�d��̠}�A��0�h!� ��3U]�Ʊ/c���'��L�@3�<i]���M��>�7�Zn���M�i����Z$Im,��2J0Qh��E�A�$ˊV�g?ir�e�Vӂ���o� ���o��\�nT�.	�������S�a#�#C���s�|��:� �A���G_��'� w���b|����	l�>k����sM����֤!��;2�Es�/}������H�׎2���ф�7��,�Y�	f��H7̔N�b<�7~�&|��:i@��� ��ćjɠ2%�HDS=U��"p��"�T�;b��-�m|]���j6T���(�q�8p5PQ�	��ZbQ�����B��"BI�pP��o�\�ށ��5���}�c|�B(�l���ؗ�7䋌�0.��������9�>Y։f��jv���eb���3HzI۝��f��2$�VſL[�~��}VRܴgΑ3�,����5�n�����҇aQl�R7��8g���o ��A�����a���t���xt!M�?s�i4�|:��))a�вf�6E�3�#t�C!�E�III���K�5<�9Q�{����3�6c��&)�BX�ʉ1�����ʡ:���R6uL��cRV�g/�"�+׳���ᗞv��S�<un�oW���SF1���/a]Q���ike�h���8[�0���ډ)pz�^O�kl��!�:�P� ���DIG��jJ�v�w���f�5��pr��Wk'�(��`�	����~��:�(���H��%j�߷�7��r�&�Yz��/E�e�Y뮷��:���CZ{���q��7爫�1��; B�p���űw÷���kY=-�Q��^;铴ױȺ��<W�$�.��m+��s��u�M$g�|{-�l�x� �%[���Uc�q�{��,���C �$?I��M�	��:�N�9���C�|��S��Ε�x+�*JY˃ �,��6���h��W��~9���2"�t�t!%�*�����ٮ�!�c�%�O������	�=�(����Qȯ��a�L��>���?Ƶ���=�̻y@��I�yhU��$��Eb+�H�Se Wշ��|fϴ/K���`���b3�4��fxϪ��^�;��X8�za�[&�tʠ3:&��?��G�e�Y��Y(��V>|w`���[a9���_���[�X�u�ph��Lѻ��'��@�Ei��m ����^�k�:{ު��.o�+��C�B=bJ���zb�9�Cy�=�}����ZX�H*)�م�Ԍ��ů���]ݽK�,Lu�VΡq�97,����E�X�d�CIU�n&TX9��c��h��/�Y��["ѩ�L�hvՋ���]!�#���N��^��<Q�[tjz�sE`8wO��Wҫe�XI˟x�|С�e�k��������>�u�⅙�2��TC.���z�һ¡�5�Le��?ϭ�V�M��B~_�>�d��tva�FYO��I'Ζ"��]7&T,8����96��h�~��MĦ��4����Ju�P�uG21�z"fSg��s�JM�f5�_���б����/����4���J������Oݢ�s�|`��l�����S��}Y��.��
ԙ	�8�S��v sP����l�L����?�}5*	�*b�rƮ4����ٿb�6ĝ�
ثE�ޱ�y߈�X��Lz0"��J�����u~x�w�۳�P�)w�4���l�{�6��!�	& �w#a4Ğ�7Oc���	�!��şO�k�̀�����ɳ����^����}5dQ����B ��?k�o���<����0x��(�m�������*�\���_�V@��I��Y��~Rri����?�gI]�ٱT�s:��}Q_�"z�9�#�}z#Ct�c�pX)B�}k���w�G0%�,)���ȩ6=�"��-q-*Wb��p�C�'�3��0@f��h�l�hp������B�2��4����U)`�2��.ģ��n��w��8}��<4��<���NW��~�U�\��.E}�������	FVc�P�Z�����d���?x�$�F���&'�D���:��a��;Ê=����GR�@�(�*�F3ۅ���T�qy�q�ӣ��Ȅ�����W����%%,Q~��������r"r����X_���FdV���n��d�fғF7����Lcv�0���{qV��*!����I����t�䍬��ucnM�;&������ؕ��9�Z���a:�sv���x��ɹ�iT��(3D_��2͖]����S9tі�n68c�&N�[�.�ފTt;B��yObd��GW7Ԕ�"��RC�Jֿ͂]�E.�#r�ª��`_�6_�8e�/���-�#`�����K��L�D���G3MJ2��B_��W�?*�B~˩�����l�Ti�(���3K���~�=�E��	u��%�C�i-W�(d���c~��ܪ	nw/B:��x�W�wW�$n��w=!� e�݈�u������,�qr��I��<�R $��כ���N�vR$t(!��	���?���?ڒ�/�wn��b����~��`�PVGm\��Dd5���Y4~�a��� /��C����N���ƨK<��;n7������7�H���#HJE	��a�
������
BF��Վ��(���l�)3C��s<�W�>�E��9W_��Ǻ�E&�*�Qw��K��]3f@�ғ=�Hj\W�۶�o�ė�p�|H�����;p'$^v��78_D&9�_԰�;kݼ��PJ��1g-����������]��=�)���g�?Ŕ P���p �c!`��ў�3�4A��k�iII�ҪBo��\�>���.��-�[IWٻ��L�G:��U���3�Ɣ�%��v#�I�P�j��*M�PD���MtQ��ni������}~;��-z��xͿ�z�i���&�<5z��4���	X{�����V�����fkz�����,P��K��kV�C�B�m9T]�Z1Xzm�7o��R#l�ʤ���ْ|���<.�/�!а����vw��U&l�v����w�t��iaS���JG�i�(�%|jY�ޱW8	̹�24�d2�\�"�2n����?P.��j�}�R�8�%��r߳����oϏ0�慩�g:�8�}-ͣTT�$�D\'٬�����C�>����&>s4�m˥B���fVM�BWO�-��o������מ�J�b�o	N��?˅kk;�.VT��S�����_\v����N�-��>���,�j�,�고o���g��:�j���W�s�>NZ�؀���-�e���>��Ip�v��"UI肕eI�T�(�$���r������^�K�ar	a�W-u�$[�����7f���u�'V������@�`�����ڲBٮ7�^���u�~$�pF��^Q�tCE