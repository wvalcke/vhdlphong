XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���⳷��û3�������\p�:�ݛt�?y6viwy�4��=�8�&��)�� P �Jd2���R{|�Pe�*�M)\�@�%�L!Rhmn�����ykH�n�@?a����M�!KmS�Av{��ܵ�l������I�,�Bp֔j��xt��U��H�(�0�#��6ftep��۷B��+p(�b��7��W��)P4|Q�o-�_3���E �;i��i��ݕ��(��~:6^�MB�^RΣE#~�����a��cD�ϟ�U0���S�� ��.|�?�h՚A ��TW��Bܭ�K�+JɆ��|�d�ݸ8|
���BN%a:���ukZ z*�� ��!fx���<�Oq����.��w�<���L~j�.����dS���k%(���SJ��"Hؔ_��6�:��GѬ�`q�tƧ�%|Z���>E��CYu8����e���DBT�ud5W�2������Q#{�8��MidY�׍:��e� ��2>ϖ�r��"�����/�ɉ&��%��E��j+|���2k�W��Z�U���8C�i%\	C��/�g4w5�k-ˑ�o�yȞ�^N;;�O;+v�3"x�C��O�yƠ	=� ��� ��2إ�v��-���� �U�\�w_@㔅�2^��!��M�n����Y�C��+�7�F���r�����u��\�_C�X8��X�J�u�M31��b�w��C�᧌+Y]"�rtW�U��"����N���V�x�f��Va�}hXlxVHYEB    1795     7b0��^2�ο���cT��j���r�vƾ��mM�5��b}�<y`�JW���0J�ۣ9T ��7~>d�:_~�.�`��K�8}�k���O!3p�a*�u�+'�M����h�2��d�l�L����J�p[�u�{?N�ޮ��Q�p��-��Jco�15Dw�z��/UJ`֚�a��#-�q\z�R8J�ජ]4��zp�n��1���h�0 ^�<��<!v���:���Y��n��w��V*ֺO�+`wB��Bv(<���wW��~�힑�|#��y*��.��-�|{�k���NԚ7�A����:�7�H$�]:-�������]�m.����<�Ͼo�J�j���n�Ddu��
'
ട�zJm��*VD��6@�F�g�"�����+����Xe���*N�W�_G/}�j7�;�+/|��lCQ�Q�+Cf:n6�zU{y��"�Q�T�30��'��O�T�ÛP�v��_zp�Rq���Xi	O-Na
�è�1�s��� lA���ZeP��ۈR�HG+�\.���A�En��H ʰ�����A��7�ș��x#A953?䵮���h��Tn"A����������n�}�l)6{�_�?7C�T`�+}q,D�[cV �������Џ����Frj
�4�Ǥ�@�<�u{�k+�МE2��_�e��aO(��u�5���3�lLd}\F�P=���*�O���"ʹ�����ɑ��cH�'�!����"���r+��g�� ��\��+��ZT��ms6�1q��%�����M����3���0�-4���Y4N]�ע<e.ֹ]�[����a�4f��j2B���W��W�sXM�fqJ:*)���=���#�63*1� ���-�<�I��c
�Z����ʧ�����H%���h��3����D�B�B4��6�>G��0^�����:)�w�m&��z0G�x�B�Uvo�'�s���*H�Q������ ��d*�h��*T�� ��E���>nM���
�Rl\c�B��9�)m��>Y��sfUi�q��`al�h��;��顊�����OY&���z��A�嚧����}xlA.��Ţdc��75e�܄�����i{��TG^��?������ȷ7�^X���К�!��_(E��sQ�PX�?{�ug��^����	���Z��:�f M��qvcp��� ˿}��������ܸ>O"�]��Ȫ�YК��Aћ�'9#�A���/2����o������_�`fq�gz����@�gd�#'���"Wٙ�7K�=����em󄄕��p���f��eST׍�F����ח?�U�r����\~H����6RC��#`N����6��[���	w/�����oB����2�g��2_�R��_�Ut	�I�%@���ދu�G+����ҭ���;��(�H�	��m:2�|����\3��j�'��0�U�ݦ_�b�L[;)�?��z����s��J�C���w�+Z' R�~o��oV�[�o�ެy��˓�=�@��� n>!��x�����nf~sQ+3�]����\�MA�g�[������������"�#���qi�Cg�п=R�Z�N�����ݐ2�K.�DtdN"��W���C4i��.�<͞L=gLr�y��f��j�|Bͱ�Il�����~�C2�a?S��'k+�	�b�.+���s���ĝ���q:9}i3�~e����q��Y�&��f���dK�y!�,�Q#���5a	�'�tn��Y�ڃ[�J���%N���c��Hg��8hdb�3t�魧^����MU.]���FNh1�'q����>*�Ƣ��}!,�����6�u9sIek`�"�@ض���R�?�l�Du�ޯl���}�6ݳ�|�q"��*��Mm'X�8�T���)�5mi�J�$�sXT��d��KT�[˼q0�C��1a�k��