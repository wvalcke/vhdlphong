XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���\�97�0[�~~�;��TU��?v!M̋�^�}\z�o9���}�ӧ�4��ˎ���u���|��,ANKs����,0��L$]�1� �i��:@�܌N�d�U�?�%�i.�	���蒼��Te{'%>
ޓ��AH�}��#�P6��/jJU���Go[�ۦ�T^(2��
����G�@�6_|K�{����I�;�I5$-�UZ��� ��`�H+g��1l��<�'(>E�_`�kE'~%�abJ��܁4O�e~�Y��Z��boi�����=����$ݷC��k���p�A�G�)��=(R�tiy#�D��p���j5,�l������²����"O}�l�:!������4���#I�>��߀�]��e�dD�d �(����r�6����p9o��	�
�ӯ�@��潵+�j��jj96����*(�L~=�Yw{sy������\��l��,��A|#��Ix������q��2aGj��~��
o��X޳&_�Xz�x�+�Og�,�?~�Ҵ�&��_�9(�Rt�G-�Y\܏�6z���}5��)�;e�0�5�R�B�:v�
�y�R�
HX������Yz>$�דp��9ѭr���k��8	�!��������u~�lHC??R�lwnǜ,�)V�b��?�h-�2ka�k�f`��R�g[Ǔ�`�ci9�n��d�pĳz��u�� ��z���m#W�"�SKe�Q�
�>7�#�X�e��0�q��O�|XlxVHYEB    6e28    1620*�����e|��u�!�������J�lQ" �-�Q&���þ�����C�C�����/5e��E�������}�:aՏM_]&������e�L���Ε"�� ����l��&srl�4���a�U���.{N���Gww��d�l����.�ƪ?�h��K�j7�wR2n�&���P涢c9��KR����#��ua�䑉�!����`��Uސ騷�0!���9��$��'�W?�y���5	��<Zf�҅�f%n��Jcp���bUPG��N�\Q�[�� e�0���f�,��E���)�J{)j��/�T�\��pj#��{����4%���K�>k���A(�a,�Y0�^*K��)���44p���^j���0��[V��B`��TT	��(����Ǡڵ��iH�\���f$�S�ƾ[C�ȹ�i�	�?��v�q�:Tq�U8az:>���7��w:���!�6�ï�Ct~��4b7n��G|9��F|��Jp�2��k�3�]ְ$�阾�C�"t�?���H��U-��_b+�Q9�=q4f��7���@�<`F�y�q�����v;��I�ZZ��(�KV�<��l��#��iK���޼.����ѕ��/C���Nim��^*fN�G/jN�	�`N��$�گ^Y�c�3 �ZQU��Q����p°&P�J��ui~�~�g�F!���N\�ci%:�M�1��Z�K�87jH_�@_�1M:<�wǫ�(!,e��������F=@dh[���Vz��փ��2�FFW)�,�		���n"Q����l����a{�V�L��K�`-�UG����:��r��&����������(rr>3�>tjސ��<��0�/�`�IL��R���W�p��s��(���1lԾn��OHrrU��Ϝt)�����Ì"�q**)��:�P6�)�[=B��8M�2�D<qg����(��fsB�T��M��qDA�����Z��N�؆�=�\�Nhٵ�<���k'�lV�u�?����&/eI���}i����s
�a_Fы��B�zս4�����<��*&?��X��J��H��6�Y���yr�����^"V�2����t����K��Dzeܛ(��JH���%�tw�Mԙ�������iIlr��;뷝P�0��h�U|��_ض��zQ\z?pN���[�"�.>̬�2�5h8��P��^��M����`�m��SXj	�7d�0�IJ�b�dr#��Djyg�-]�zNpt76�׿h�h�R��U�:1��~A�/<�S�1��,8[GuCq�4�y���c��0W���L`�h� ��7	i��ŉAe+��FR��Aۑ��u�f�]�.�b���LҦߺl��݁7��˸3�ݼZc�{4I�W�0���A���(Z;�w�:��3��*�ހF���9rv10]�m��oG��Il.2����M�����x2~z��ռ�m%I�By���a������c� f�ݺ�FKǛ:�kt�O��:YI��kr�f�G�������evw�� �+E,֠c�h�2H�����;.%�ִد���-���"�k���^����E��}�.=2lCV��O亝qsr���ϰzb����,g#�іH�X�����MV1��e�N�����e,��s����qi?5���C9�2J'3z�KPR$�g�j�|ԣ�fB�$�����ވ@f�!3s���͙������6����>���ؘ6��BU������� xb�&x�M(�	nܹ�<}s�Nҥ��;=W���{tʣo�	E��H@\�l�k�m�Ք��-��R����Η)�2�ڥMf,i¿������U	�(O_�ZB�oN�餀�v2��5������~#Z�u&�3"NIi}��WΙֳ	��}"���&
�����\7/6�.�I�3������0��c ��H��dF�"귙kJm�c�<ެ��!�䎔Ò��u_�E���U��P�_@S����� ��4@���e�7P�X���T0�@I�?�v ��a�V���C�Ng�&��2py`8����+\j_����3j"�߆*��=��*F�e%�c��S�~Tt�ZGW�k�ǣ9A&���@��'�zGA�R��0R�!�3*�%Q`���������n�=p����'��>#��2�O����zq{�=��2S�}a�� �d}W��`C@V����c�[�|?��<G��-O�����P#J4����*D�O����b��e3�:����Q�[�	1�ߕ+?�p�ew0v��}�*��!J����ep$@�����0~Ư��:#�-�f���P����CC/9e���"���Rs�Kπx{��`Дw}��pG;! q�p�����o��N���&�p�,�6��p&�cǷ*7��r/�L�� ��(�a���.z$��ss����?�06�1���(��?��Ŏ(6�d��2^��TF�M���$-2����n����IY�nq��WМ���C��o�)c�0��h�E�i��Ȕ�D6����6-�J� .�B�rI�>�|��
T�t�_��#��k��:�'(�/�Q �3$�+��黎��L��Rx�ÿ`8�w~W�қ��CX�y3mQ�������,����%�M'�9R��46J�$iEF��1�~t6`������i�]��3/��/�w�~e0n��|Q ��Y%)�m�)����'dK��{/ھ���=�j��L,�e��FZ�	� ����Y@6�`�����(���U_�����o��p��:A~���Y�H/���Ӿ���t1�O%�J3m�>°�o�%��h,Q�w_�}=`oI'�R?�f밚�G��dTs���jx��>Ef�u<�4�MP�O��7~{��h�OY+�d���n�\-�{��>���
�i���Գ�H�0W��s<S3j�k��'�����/�}��}/�y��Xf�9�Q;���v�J6i�MN$�b@`�?�����,�������	� P/�9W�2�'^��V�e�_��e����=�߳�{�#=�(��}{`t�lW����(�I�� Su�9��d�|�qA���xݳ3\)26d�����:Ţ��|�9����i�Z#
$���ٮ���J�ܖ�`���� ̆G��]��bB*&�Z
�ʛ�Jt�ׇ���`V��~gP ��bs��Tʽ���ZFұ{��Zv{I�t&�9O8��d��ms���7�w���uėJGTq{t����*�w�
h�#�)�&�����ٽ�Ǹ�h 	LѴK�D\�!�4VTcI��c�X�PԬ�I��k���O����>�rt� V�����N݋�;Vm��3�}�q��F�jC��`?:٥��� ���iv�V�O'�e���Ӊ{a�@�J.�(��`�8\׉h?r�N�v�*�4�5쾣]����?����e�jcoB\���ᐓ��T�qn썘0�0�N�Ґ��yJ���7�b���&�{�CCh���^%�.�߂���G_�k����9�<��r���}�R������V�mu��=7�2����	܁�݌�S���P�b�q���8}��������Ut�Dr�'e�x�5Z�8L��zS�����,��φnm��� �|À�m�J�o;c\Rw43t�һ�k�Ṯڢ�`��3�9N%Ui�	^R�y�, - �J���XR#�g󶐗�QC����_x�+�D�ef�����|W�֝6GF쐪�Qy���ɫ;(�
C� -�2r5�WX�R�H8�y�\��f��n�\�K� �S��,cjώ�_�z���:�E�m|�y�P	����$��~�X�M�����.ށ��չ!�q߷���.7_B�@�V�?����U;C��H��.8�8�g������ƊB�u$Z*=��V��v�@v���.#[<Qq�'�{˟��bʌ*D�Ϋ?Q���z�yW�?$��W;v��o��VI�/P!c�6�'tԏ����U8�ja���C(�@�:g���S��'�^ D�߲U�t��ǔ) �~��n�<D��n S�b��{��Z�� �@e�:o)"��Mv��.]��m@����7ĎLM����r���5W�����ds��*[Iq,�-��i_r�jQ��(���Ğ��!���Ϭ�����z�?QLc�XX�S1ԥ��/GS�Ȣſ��]�zo-�i�\�T�q��)~�Bf�Q@��%|-FCCn����eVś*�T ݊#;�H�.3<��Q�y�����L(��i������0�
�����+jߥ�e"t�W�s�#X�df\�~0���֑� �E=�.����U��NI?Q����M�R��vB�\���Z�k�/4�/F���$��e�����G{e�S1;0	�y����i�fn{ɲ����K��wT6�s_����{@2�6�.+U�iZ/��T"�%�q&�\`�+_e}<$`���'����0C[c�{,q�o/��fE�ڵL�u�aM��� ���n����Y���7�g��t�S��qU9sG�Z�v��[6���f �;M�'_��7R}�W3i>Y"��hepj�:��Q{Y�hs��6>��j�R �::B7�L(�yDo�埼�������.`b]U�P��g�.��9��纹%�O}�g�xE�"�ק6�<^.9��c����1�Jfz��'3�sp2�Y�Q[�P���^����*>����	�;�bB9��\��+*����Σ���Bo�K)Is��[hO�94W�J��so��$/����D��\��K��2��㊄�� $6A@��B �ZV���(�UQ��`)*�m�ZC袹�j��CҴY���*�a��s��������♘����ys)���ok���{MPI����};������
��|=��`��# )�8O��mrAtD�����^q��-�-i���=��{����w1*�X0#���)@G��v�Y�F�觟�����˹�C�j�6�)R�fx��f�"�չܓ�e�+��*�l�-�����TBL�T8VqM� b�%�rt�����b���R�S�.���ta��<>�s�t�LV���@b����H�"�Ǩ(�t-͊��z�ڕ��X�Dׁ^�=�P	p*�Т������$��i�@D� ����la�d���	W!+�w)��Za����H�p
YmF��6��ON˴_���4���n���6ѵ����5w���o�%����S�����Ɣ۷���u���lo1Mm�A�@��T�!���-|��Sl ��yP,�/����ɋ�B���'�IBJ��2#Fv������.�Fk�@	h���
�����yڎ�Z4e엘�=sY�^ޥ�"d���!`uN�V���_�p������=#ǰ���7��%��F��Y�C�)���mў�9E�|m�Il�8���]	A� Rt� �Rf�[p	�~��k�x75���� �9���q˨To�JS$ZO��),*���70�M	YCϪ��ҵ���rZ�5��H%�?����N��?�:�Ł��;��ԗe�u�'��0��]� n�E��̗��Ŕ������Ϊ6�uU��ߚ�'�E�����8�w��"�vH8