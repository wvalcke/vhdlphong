XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���~������V684�QHz�ra&��i��`\s��P��wJ$���,~tO�ĸ�����DG�9߭>k�$ي)�&Ԝ�مtW�Ow���{���7߹�l�q��k7������ �(��?�Y=� n����Y*���^�2�Ad��u����XM��z��ņx�t6�vJg�YK3���յ��W�� _H^��8�&��Qs�{��L��:I��&v�����e�.g�]?Ӯ>�7�|��:䇎_���d�d\4]��n���9��ME��*���T��J��7$��!.&�e�^*�ŕ.�'´h�Ѥ�d��F]����w��p�g���Q���j��x��� �\"��",�Ӿd�[�m���;���o��Pm1�Ԝ7��-S��O�m#���1/wpR>[�<��>�զ�k'l�Οp���\�mI,#���G��w��<�&)�M�n{�ы�.Om���1-�}����m�ch������vłК�DD3" u�&����Ĕ�ۅ"�M���Kӧ�1g�PO�J�!�����T25^�a^6$�t��ס_��g�ڌ��*h�M�ٖ@��i�9���}1w�%��b7r�� i������_)-��4g�j�<�w���? r�3����]�2���x���p,H2,��X�faa�#e<��˅��iQ7�??�`(yˣ������?	IǍ�
P�O�ݻ�$���(�d��N+��Om�N팰�͖�Մ�w�%4�����XlxVHYEB    1602     7a0C9�2!5�`?�Ġ�vc��r�B	���_�����M�a�cR�Dq>ݑ��+���(3��Bt��V'g��xd���1i�����e^���5����-����[2���W_��ЍAG��þ��P�Tk2����7���u��W���>��p�Z���,:�37Ԯ�ݎ!=�A��tU0rm�Ep+p��Թ}�����x�2��`��_��EQz�y�啮EHu�����ke(�g�(��u]�tFRs�7�B���M
w�s���i�euh�Oߜۈ����S$o ��q�f���E�e�bS ���>��M�&o��������/�2[6N9(+��\��z�Z&!C{��Ơ��U
�o�U�C͙:�D$����z�K����)�=�&[�l^����j������O���L���q��83�}م���&�WVѮRB��&L ��g#3��#~�!D�]m��#�sY��$vSUx����H:م'�$���&��
��x�~��gk�����p��#,μ~�:�E�V��=���9;�$H��|a�����T�R�zH�`D�Ќ���?��}�݇)8�[q�->�J�Z�:�S�>���|��Xz��mD��ʽۊ�_�]z��1s�����biw�KT��G` +@�*��[0�"�2�9�p@�x(u4��Y��~��3�����%�~��^kC�rS�U���&���Sm�`#X �	������G�;�{��V�F�Нv���ê�8g|ʶ�z�<mU�*-�}��{Y-���fv-F�U��Ͷ��+���Jq�G��kj{%H/"H�i�9?#�Ŕ�%����R{uC��3��&s����9U#�Z��v�f���^ �G����H@c��W �(Á��`:��4�Y�?��*hk���A��.����3�N�mH��B-�SP�����C�eڀ�zz��U+�%��(�*���R���t];7�I��@6d�\�N�%�:7�K�I������M!n&���D�oA�����G{|�#�2��A+���i�'>_���!��䌭�k��y�_s�V}�J����։�T��ۼ8�4bZ>ƻ.>*���r�R��\��S��D�YI��%9�L��e��e5�X�7�{=���B��|�(�?/?x�A�.P��9�+��)�ظ������6}�T�	YA���?�1��ߕY�g���Kwc�.M�4�l6����G�%�Q�%����z�����7��l�R��5���`_����(�L�6������l~*P)t �G�ތ����}�����±��2�c�zɑ� ��ya��*�l�U��4��ϫ�կj�F���)�)!��E96�3�7���|D�{���ŕ��Į`��wPd}�\�U��y����ͫ���׳��/��Hx=赐��M�Ȟ�%�� �eI�2��@�#ڜLD$�4*=�U�� pY��<�>j��Q$ѶŦ���<:��J�@=��V�.�ܼ���9����7I�gM�n�	�F�_���E��ʏ�hR&~B���Sfd�I����D��K�)��WLI�6��,��[�vg��d��R���2�wz�6�?껷��6�%&<w�0����i��>���Fd1���L8�g�W�`��0�|����C�螒�26<`'��\ZN�+~%��<&�F8(1H��:��%8S��ܷJ�E�؂a�W��U�O��3ʹ��w��*��#C����C�gM��V=er���>q��W�@�	�����/ԩ�3Ⅳ���������,@���o�QRs��S����w_u7�����yJ1���sUC�K��	���F����ᾏ߿�ݣs��<��W�ϣ�
�ұ�P/%���޽�͒�uG�g?���r��>DV%�7m���&��zP.��z�����qO,G���#�,�!����j{KQSb�~\_��VpZo