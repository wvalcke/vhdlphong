XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���>���(����ks�	I/tR7b&���fR�Q��%d� k|��D�L ���Eɂt�M��N�;R�l�B���0<�v���]��}p͏��*�1�Qm[R�뤆8����e��; �wĬ�J��m>z�*��8��X��Ĕ��W������(_�����E��&�脉�,���	��a�J�}����P5�s�fi�]��
-@�-��r��6���^VC��QF����Rd�}=4L����=�{�{2:aO��7[��H+�¨�F�S���y�n�T�D��G���؀����5��c*W�	]��%�ob/d:�qOoO�t��)��}��W����FC��S�t��f�ku��q��Ӊ����&O`#����P�r�,c���7�u�ç�o�v�w0)�ֳa����ب� ���U�5��JX����]���3���G��6Da���/W�sbi��G��(1�{9e�4h^qV�d��h�B�Mɑ��x��w������>K��n��jv�|D�hD�P�7$h��xF�{���H���2�C&�+�y��\X�(��ו�?��tL�=�\h'[���b��	�$���1�ƕ0�������f���e�7	-�pQQ%U!H���qÌ#����䯶a*��F�_�tK��E����ǣu���v������^E �ņ/b��'�	�՛�B?IV��9��A�! $"���&�%X~��G��*�"��)���1���.�m-p� Vu�RggH0顬I��fXlxVHYEB    4ba0    1230lM�/��~�H���r����Д��2�"PyԢ���Q޿�U~����;�i�U�Q��ᥜ�ؤ��FS@��ȍî�xQ�v㩯j%�e8�P<��a�J������cm<�d��?��	A�AkBX��V?N��hc~dH��H�/��l=�5���Ҹ�̊Sk-�o	0�+��9�NIh늽�aТI������&�^PO��vD�:��F>G�����	Լ�m.O�AG�@��,�n�A��!������?�Zy?s�ĸf��0��<��G��c4tezbR[�E�L$��!�Q[�B�~N��� ^X�M���0�p����f�,��9P��lQ��t5�J�H�Q����+�q�~!B.'��!a�;�|>0�d�-Lh�+��&s�����1��N�r�ӞS�OA<�&����5��y8�<��!�׾!�}J2�4ɖ �e"��{*MrQ�u�溂��������&^�@����_�0t�eFRi
���7�>!h�(�-{�l����?�YJ�.��%1 �P=;��S�W�ꬌF�����������6�(����t�^��;ԖԔ��B���YK�v�P���m��0��N	���J�c*�dlj���(L9���PУb�E?{Ė�F	,����MǏߜ *^��r�e���{�����^��m�e/wp�t!�s�g=z�nî
�K'Ig,v3���d������~�n�>��x����tE/���Pȋ�/dL�s����>��B��B�)">PuI��G-A|�2�}������U/'��}���8F&�����j�ː��c ���w���{��4�CV�Jk	����x�/��C��7��?m����Q�=�_׾ɥ��6���<T	`�S6 x��t8�(*	�a�!sV����ґĲZ�$�=t�n�B�ɣ�
��wf�\�ix��������%�������ĉ?��H�M���j���f�{���.�ti���ʟ�89���5j����ģ����⸥����ʛK��jz��)Ċ9�����.,��iX�G�ʓ.��������&4��F���Ѝw�>��5�_Mqg裈�D��BD�D���f�?wƷ �?�)�4�?�Q�o^�u���07�Fj�Di0���rhJ��N!�z�%�&"B"��;X��Ā�±�"����*!����N��5f��xs���8�(���șt5#t���9va�%,��w��"��K �'��x��Y{(B%�H��L+����U4vu zO�s=�U��}�*-FU`aw�H�B�6ڿ���{=�)�!b�J��Q+Ơ�'-t���{W�y� .�J�,:�����ݷ��Y�n��I�2�ޖ�J���J�Ei��ď��.��Shʁ�����@/W�$ϲ���M��ʉ<@D��$,�{]t0�}ߦ���6Q
!tH�-�[�E5#jS�ą���Nx��4e����y�Ѧ*�`����4�z9X�������۪w��2Bm���=ҩ͛/�K���k�}�e@i��[@Γ��>4xh��PkK�NnM�<S����+(�KuA����*�Υ����wq@:{����h����4:�D�I���Q�|鈮���jU��s��+�J��H`34R�vމ�����4�f�bi8Y%m�.��i7?n�:���r�V5����|��b��WD�LݢDB����Y��@V���R7���X��Ѷv>��J߀:�ӥV�&&�(�Q%��GKGr�l8u[�x�<���~���#`�F�~x�g���*��erLrb���yݺ(��M0˔!%��+��
��ic��1�Uu�0�v6�x=f��d� �����6HgE��Iى��h�4���q��b�4Y;�Zm�8�4�,NQ'�
��N�L�;�}W�\5��'=P���2n���l��x*4���#� �+"��M�'��� �Z�.P���A�g
�k5����i���4̃u)�yy� ��9��A'�X�~\qۚk�{HA����Ѣ���-�x�VYr�qn(�D/�,:)���FĹ��܃/�X��"������d� ��oq�E�wf���i��'�CqNP���	�J�kn��XD���cK�����ba~r�o�'�:�XT��o���p�VZ����r��\�R���Ke�����#��Kc8�vJI�Zڔ d���>f����^�T�?z�_wj�#�*G0Z�|m�dM���:��
�� ��kAK�QΜf?��ow���XO����}�nl��ط�P�՟̗G���\)�YK!`����v�C�/Z��(#pb����fi�,��Ϊn���T�GǷ�BCk�LU�J�^�T-N�
�cj �8���0�tS٭�)��XZ�m)��ȡ9���U{�����Cg�춨-?�J#W�O�1��A酊�X���{�wF�/�%�y0�,���S��G�V N�'۬���,��w{�%�\<�@�4zk����?�k#�0�s�dm��/c�O�r�_�»[�-{Y�*f�����܁���(� *[z^G�W�o�A`��(�M�`/�SͤO�0�?�-�t��00���"�==RlY�]G�\3�ш�#Øyg�k�u	��_��k�@B�w6in~W����oƥU�0�}ΰ����N��������=�ʱv�Ľ�Xq�H�\!����~!ΩX8���HX�(����m}�+�[pB� T��B;��� .�_m�
�o%���ҭ@S2��᠕	�	�h;!Ffv����<]c54ӓ}���-n`����>��p@�n��������&w���c�?5a����Z\cM���tn�!����d6����v�tO�m�/"m����a�;�.+Yj���u^����Q(c���7W��\�nj#���͒��x�:蜶?���!��L�471%��s�G�M�z��{Y�]!Z�#�1Vplk�X�m����ȢLw�/��Ճ.�CcSuK�ƬZ/�SU�5Q�
t"����Ii`�K����U|�E*�s�@����oF挪�c@q����>��T��W}�">t��M���+�zy�%_�@�e@��s�5�P���U�}�����Q4�,�޿����������M�Fd��@����f�}s+�{���ܐ&�UQ[��uY�t�(��y��0�G�x!gR`<beφZlR��K+Ug���`�䙂��\�۽RǱ�>��δ{GM�=���J�K��mb�wO@,�睌�s��t�'V0����8�8�*�a�H�����P�\^���D�&��������2�����{�2~�iִSƾDN"ߌq4��wUq���œw>������Ҕ��[e�;��BX����z�E�	��\�i�C�~�/q���g�9��U�W�E�;K^������D�详���.1I�S�Z���9;����מl�Ƽ��熘۾8O�u;v��؉���׉����L�<sI��������4�B�~s���˵�^���^�~-
�l~�!h���m3�.�ys� ��$����b���8��ʺ�,�v
+�W�8Ʈ�n�3����:a���u���n�� O袖I�+r== {�%�ף+���`Xa���)��·�w�m7V����d
�����('�>ݫ $�����.^�E��Ͳ����4�Q�J�+`pRP�s�P�U�%�"ߨ�	ee���Qkd�ѭ��"4+��UE�[�����,��Ͻx=�d�UK��`,�U>ph���Y
���ĸ��}}U�%���:��_/t�?0��*ة=�Zĸ5�:��w
&\�1^DԯSVH]Up�/.���r�X����I���G�|*f�bo��<��?V� �y�S[���R]�ڹ��$�3)��7�R��˺��8�E�X�k�`,Y ��5\�g����[�SV�)�?Wn�
��6�O���D��a����\YL�Ew8�@Q\�H�ˑ��������V��)����,�.���+�3�m��3��r��=�Ph��-�}jpÞ�ߒ�D�/U��6������YXL����N�'�YU8�癕���.U�����ר7۶�\N����Ÿ��2}����2�П�r�-|��g�mn-[l�����;����g��\����M1���w���
��<��T�o�Ѥ�	4d�,WOF}[����=2V(�^�%P�ȄPF����d�� �hN��%��;��mCh#|�{�-7@zCii4�#��"<��.p��ZFJ1~����V[��=}h�v�F���tE<-��sB" ߈�#�4:@�^�_Ǫʫ.�V]��@�§����~��K�<�1��������1��T+�U7�Xv���BK�����݈}�2��a$+�����s���?�ٿ ���ܾ3��Y�D�BC� xk;lN�@_v��U��d��������sW�A+�|�mTu/�-x>X��DLgȧ�J)�g0V=8�6�b�/ ��k�oΑ��o/������;�[h��ꒌ�<�{'`,������O>�y��{˴��î�YQGr�_���rr�~oI�VbU���t��K��ps�.Y�S�8U���ef69���u��$�LX�