XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��&CM����"���6����!d��;d���rJ�cYi����o-����^�;��s�u4+:fո0`F�6��=��n�U A�!��cyH��~���ΰ���ZكSY�}�i��RR ��Ю�Üs!�6���&I��y��2|�O�\lZr��0*,�n�}At��{��	�RO�Rg��J�{�Z��z�=Zo�@'N��0� �yo��P��z+�L�2�}��d��cڑ�?�`�{��0�X��S��uJ��K�����W�G�UT��d?w�Y^�����W:k���D�Fv����/c�f�1�Cݽ��k5�����%4j�In�HUe�������ә���d���g2��8�!�Т:�Y%a=����(����
����x����O��l�^e�pt��#K,�*m�&���ƥe�ݮ���:e� ���$jc<���=�zr�f�K�Xp�$������F]��U3��j�Zo�w��^V�8J�7�ݔ�*�M4�OQL7M���}~-�M�2"����a6Xt�s1V  [��H�tb����X���sг{04J�-��Q�i��[� 왾�ȾspP�(`�$JN�T���x�_��Y���-�kT�$z�X�0�Gb}6��I5���9�#��;/A�jFiGZ�aZC�P�7�������Dv�I��/V�|MV�������[1-�K�#Cˢ�+G��
���Ԏ��Z˘�g�f��;�}�U��&�&��_�B�$f(�УXlxVHYEB    5ee8    14d0� ÐQ�_j�g�l��{�>0�*�"0�ud���0�H�-ȃ�<�8��M�_����}i4zV�M�!e(��K����E;$���zU����j���-�ዧAfnQ_j��|{��rm�:4��o��ۋf驢��z!��I`gCT@�!GD�L���͗�O!�c���I~j��O�n��\��h�P��.y�L�U]ۂj�8`�~οT[������m";V�� t���I��2��M��cp�;�NI�;���o��$*�x��W�vUG ��ڭ@�x*����7S��RZ#?B5�(�w7��cV� �iU�h ��X+��ק�m_j��?Y��O1������޹��w�n6Àݜ���(9z�2� ؖZ�$�2����D���&i\5vN>�u�Z�,�m�L�T����!`�O�u�|j4c�O�����.��D�b*T���1� ��-���q��q���Fc�;nK��sQBc/<)��0����&�
���Q��/o�_&�/�Ծ>"�\��f�w�T
�c�ej;�|��o�8����I4���Jc��g#��Y9�3+d�}��}���7哟�Mʿk.2��m�r �_�x��a8�8��_qL|�Rꇜ�1j���"lDf����n���r=�-hHH  ��[�`����M���P��k����h�¼����""ˆ��4��	u�� ��/`, �N(L`I�Y��Ga�u��&��9|'8x�E�䃉n/��G�de��.��V��`�mz���+;�U��B��k��6St M����w��������r�d�e���<�%#�<�ʉ�Q;���ԕ��n�����*D����9�Ak��q�^�U�gND�D�� ^4GWAt����C����a�),��K75���'S�@��4>��V�{����2t�$iu�6l3���o�\��)$E����JV��zF���o���9���Z;��]���L�ҰpC�ۄ�	s/���X#KZ�D��O?��C��uJ��)��@}LrS$�~|l�� U4I4jAG���SCZ&4>�$%I�[ёQի��3>�2�tCnq��|K��XCb8`ᯔʢNv�n�u��"��1n��DC	;��k��5#���'��'R}�y"����˷|}�^�s�3N��O��X�]��5��(��^Q��g! 	p� �������s*Y����'�}�賧@Yz~X>=Y:\��A_>;�KsSI��^/�7;Ø( r�c�H��~��⏱�`����$2����xB�p�KB3�Na��y3a�~H��B:�v�?]������t�zPb�h 8Mŵ�@j�`�}nq9�Y�E�׉�n y/��"���C�
��G�s�s��#�pB�66��v�BT,�4����}k�ǡ��貜��`�µ��g�=�����V�6TC�kp�lfVs>��~q�sϻ������J/*�\!����]�-q��q�������+��ݠ��Oa)�S��c����/ޔ\���3s{l�f�8���!L�E�^�O�1l҇�:���$�5[=�����v���B� E��]���ۤ��S�:�PFb��Xc����)�gG���>�N��		ݪm�Iz��B�6n,k��˭h��oK�L��y�4L mK�ݜ4�n^��ե8 fiB�5�q�����7�ɖ:��p�/�D���6��*\�ͮ���������3�nuړ>Y{%�R;#L0 B�ը��B�ڛrQA龹N��n���7P�Β�jlz���'L��ѭx�H�����9��Ğ����M�
�Sg*b-��%��Y{�oȣ�p�	�)���\���DW9�UKj���1��,�.0[��9t�͎k�ڠ�����g���"��J�Ь/��)7��d�Vϟ��i�=�-�Sq�7zY�\f������-oD�S�(v�26�O}9�2����|͑�:D#�����T�=jq��T�`�������3б���Ed�5�c��b�����T��+1�����j}�1%0�٩.&�]lu"�==n���ͪ�A�ؚ�sD_ˊ�X1�Ձ?�ï�D���%&4��.�	n�p{N+��-:�.���)���-v��ga�H;�L;n@�a�wF��|��ӎ�E�Ha/��Q��MkG-\���k��.��罄��.��TY�Z�$��Q�0�7�X�#6y���C����%ώ	GU��PnUI=+(�Q�zb�u�>��H8�@��Rp�]���t�B<�ƇH�N����v���3������!��<>�_H�)E(Sg�~�x_���2�S���I݌P�p(�^���l�+�^Í����Z٨vNv��u��C�)��rX�m@w�*[��U�n�� t�����"�&��bڻ�$c�cv
B����L��V���켑O�o&�Av�����8qި�6	����3K�F�窫SR2���<H�:IQv5>�8��1�g�q6�
L)`�N2�4�����f�H����lI�v��oK�= �n�+�?�8@���M��0 �� �o
�F_?�99Vj��)�*I��(�[i7`�m:aw����tȑ,��_�D�!�$� ��D{}߻�?�[��OW�R��,��g�J���b�"�_�����j&�P�+�G�+/��P���b�)�Ĵ�N���ȼ��{@�2XX!7U^e��af5,&\�}��q�
Dk��
��$dX�^ل1����'�'lI��Lu���:F*S%:p|��1u\��0Qu6��D�sBnR!)J%��9�4�9��WY6H��9�9ӡ������v�$ 0fT����fs���4`I����h���ق�u�?�u����C�JU?����Ffd&չh��%�\�L�j�'F߭�����Q�%�r\	��"_ߠb�v�73>w'�Pax|�2)VS�?L'��ғ��"�)����-�`ʂZ7���8�[S�������k�`5"{.Z2�A���V�+��/�{)N
��Q�~�B���n������_�g\��Ga��֖&����u�1a5�pR?Vz�ڬc$r(X�]6��y��^g+�f.Zq�e���{N��</s�?Jn�]�N�v�`���8�]��hQ�x���_ոY&�u`� PZ���h�,��Ѡ8�k��+P���vg���3u ��ۡ��Ә�=�	��S�t��`f�����y
���F��a<��k>`H�ܛ�+�w�<�T%�,��.�����6�����;	�%�"�:�1°A�@ϲ��I@5�;	W���׌��X�E������o��ku��L<b�b*�8��B/�\������v(]ϼ�����0n���N�	�"y��|6�u�! ����T���]W\�H�/��xj@���CR�U,�8=W�u8��\:*���/�t��I��_��
�C��G$(ذ+zP�ɗ�c�8��:�>��l}d >�M-���ڭ.E�����^k�lO��_ӺQB�FT�u��emg��7q���XW�g>�-�L47�;�Z��2��ρ`M�΢w.^���U`���z�T��u�L�n����C�$x|�Ӥ��h|�(�Z�ђ�ȃ�Q s�d ?��/j|[��`���̧$Ȧ�;�������%��Q��A�����|�[,����W����u���G!$K��ɷ=���4h��!\��\	'��C�2S&8��!3i�+���0ռYV~9^������_�1G)5踛��R��2,��w�c�}��,ǜ��f�tq�bלnU���O��=֢$u��	'Ȥpi<Wb��0��P�d�G�l��9Q�9�2�((�!V�x`^&��l�
&d�9C��T�nN�٨Jd�p�y!����GעV$�Gַ���,k���<��{G�cC?ӗ���1�N�ʌ��»����^��3E6���qm	"��Bgb�R~�R?�Q�K.T�4B<�K�z�2�fBK$R�]ж�|��p�Z���i�a��4�~����̅S(��>a?qUq�������s{jet[��ٶ`�R���6Xݷשx��F>�Tvܳΰ'�z��
?�Aܻ��J´�`0̸y�$������v�Q�o��>�P��x����7���ik�{�\m&�]��|�"� ��	z�#��?�2,�2��R�{t0�F����pN1���j�cۨ0�g�3�� ��>D��ռ�߂F�M�����r�7Ǯ�r�0�Q��yh>��ԏG.�&"X�����0���*d��=����d�o�"3��-����GڂH�����@�������/�ٕF&Z	�a=�
�c�H��[ӿW�D'ڢ�G"˪��3��4\�u������)+D-=����}e�\g�	Y" ҏe�x+�)r���Kk������g�zf:�}�Z��5G�{ u"ɱJ�)S�d�l��M�����/��  ��-�d��Oɭ��g}G6�l
X_Y���:mC��_�<}�����@k�A4h�:���H<�=$�$\�#���h�����(��ϰq�q���8�����b��gض�N��|�H�l7��[M=(�'ɢ钵ȁ����MD1�xT��ƗD�&����N��%�����q<�^��}�-����>kK��
q��-0VU7�I�־�/���o�����3oU���H����!�u���KK���w���eg%�TC��_\x��� z�*X��V���\���5���Fް��[�!��cU�ڸ(;���P��+>��4�߃ؚjH!�d]��I��И�X����kuR��-'�3��g̐�Y��H%��4N�͒z��`"�=�y� �0!U^GH�f�n�>��Q;$�K�a+�_�� �(v:�JjbY��&�q��,5C���-��j�@����ui�rc��n;uIɽ���˱��[����{�ڒƖfߙ��g,�˓mu��?�rg#;y�\�l=�]Oʂ�d���1�=<8Y� ����3&�w��~F;�c �l���A�="��HƖ\l�2&�p�]����0`�8=>�4�4��dn֛�XZn�u�3��m�@���l�d=����rIoVt$~�G�VCJ/��yG�f��ʁof$;�xH��qϳ�}��$�:ZrZ�4y�������Xe�I�aKU '�2�}$l|D4��$�MϏ ��W����];%�YPڥ�?M�%���ȍ�ʏ��]��2�M�9�����H	�� ���~�VXr%nr޹�Z
캳�Z��6