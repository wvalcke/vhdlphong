XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��d} .l6Q�%d��)�Šn/c���b$c$�^-Sw�R�I���#��<D��t"1^���C�'�NRО**֠M�{���l���>TdJ�R*�
��$�~�|�Z~�U�!�pJ�KA�5A�Q���4M�l���m�[7�p�sg��f�-���"��'b���A��݁HZt�nV~m���(�W��s�Y���T�̑%[�q,���4�W��<l��>�Դ�ʾ���w��0u�2�k�<0����ą3�K��lr�����ΉU���S>���=ݥ��>.o�����\��Os��ݴ���A���5t���2ɿD�Z��2�m�����`�i��1�U
�"v;M$jp���
\�0m�b�����|n��z��S�
_�AU!��t��:�~�t��h4��Ϊ��S���%Q.!;YU�<�������&K%(��ڂd�;Q�[�Xp�Ѳ�*[��.+`��u-�E&�N�
<�̱�
p�p���z����|���7�-/8
�mԏ�V�v�J�����$gӗ��A6&@�d�A:=͑�/=��O���aj�:��q!2�� ���^懻����uwX 	��N^���J����G4�۽J$���G975�kM�4�(y��O}T��\Ȃ�5����M����[�I��K]�~>�qB��=�k� ���`���\�@��@�����K�G�''4�t���
�beS��Qj��Ȯ�=���n�)���aH��m=��,8�_4q 
�\RZXlxVHYEB    3d5b    11c01E<�1W-j����ӄU���۴�n@J:�V��g�m��� .:yF��Q��v՜��'n΃������彙3|�
����XH^�j��f\ga�X�T�x���	�8��$�=b΁��΂��SB]�L�k���y�׵.H����:Y��E�d����Ta��?�`䌧&̟Pcs�8}ZsͶ ���.�p���&G��6+��6�8ֺ�sd�o�'ǽ]�-��QԆ"Q�[�������ąũgQԛ���f7���"�X��.�R��q�,�>�K%8p�C� �˭sk���О��o¤U����O�j!X�����{� �U���8���η���8	���"�=K���M��?� �	����f/��QV@���l�{ �cKo?^�X �Ě3I�(&&�KZ̳ݩ"��x��2Y!��+��'�-���^�Q����5��Fv�q�-�?[en��Cx������C���O{-�it���)t�s 8>3��y�uX,�j��mN"������Mz���vA���4�WN���)�� N	�W���gV�����r�9/��u֐��8��յ,�̷"�����W�B�i�ΰ`k�M��|X��T_v7��״/��E�=	+!�&k�Cʨ���
`n�t;��g�T$$iF1�sz	�5%Jš�Ĭ����Ag˕�f��8�&��<�"�?��a]�IqVJ�ܦ�ıW���b���!��z୲P� 1P�"�t(�)�Pr��H$,���W3WmunU�u����O&sGߑ��O!� j\�UK����'q���vSY=p$-�^�v7$����ֲdX!�C7�u��N]ۯ���\�L�
ӧ��BY`m�d]��t	)o��W��&��Yz�=7~��� ��Ǳm'.��l��ܰ�r TE�&mf�Xd	HLP��05n@kK�$�@��K:�Hd	����E�J�P{��]�~�����x	�~A��`�arDU���<�]�fݹ�U�ԁL����s�,�m%ca����ҡzgU�� О#�zRuٰJ����GV@�(.	$�����0P G7l�	�;�b����U@���2�'bh�f࠹�yvY:���<�ܟ�Z|�����sM"��K���LUN|U�;��n�ľ���i��{�U�W�\�q���adY�?/2���ɠ�E�I��؞����O}Sō�p��G0�wlU�I_�<]�e��c���9��Bo��n����(sf���_��������Z)�Or�'bF^����R2u���=�h/�(�ds1V��f:��U�m�Q�5��m�J8���!4=-�Ǭek�J�Ql12��֕���v)�*��jm�0�����1l��w����}���_m�=x���&�II��J��&��5�fP��Eb����.z"��F�q�4��t�%�A-�^Z[����_2^!�ԨL�[��듨�}e���{�=]]�יI����hx��f����)����ʦq�I>��j��̔-����Ҵ�l[��ɻ��A��Q5����j|	���Ӌ�M1l��rW�rݘkP���|,ʪ�Z���m�C�Rj��2<E�v쟭Y�o�Ϥ���]]D�,��O�<pp�/����h���/�`����5$D)I�ou��4��9�*A���Se�8w:���?�S�N���D�
\ML�t����lny�G��������8T��N���za�;tY¥ �<����:����A,ɧԌ�ۨ?��bGI��%�����J'3�X.� 'N�Ƌ�g�Eg�(&��}����4 YP�F�1Tp�BA�S:��1��Z�omYp���ʤ9y���><�bz��̄{/�ǰ�J�/D�������ы���A #	���
vH��z���)�����h���g�*[d�_���-,�ok�g�/	b0p�Qw�l��@̈�%�Ĥ9���L��26bi����3,:���������'/�Pg;���Є�S����`J�����}g��;G��#φF��3�Y��6���5��4_7B�U�̪F\��8��Tj_��%��x3_�Ad����[��V1m$��T��K/.�Ҋ���GdF������i�U���^�2�V>7U����	<W�E9�X��"[>U�UOH�CN.
�Ǚn�Q]�>�-R�p�?��oE�a�b��|����GU�G�w����+�~��t�:����c���d���𕊿qG��Z�4u�aa��މ�G����C�\�D�Ki{��iS�$�~�`�.0չ!/y�)]_8��|PM_��w�
��^�fQ��4�g�ƞ#�hV�U���Z��D�ôNB��;bP�"].]��?�//8�BA"���R�g��V��3Lh/�K���~&�kŦ�<�]+�a��NK��W�+�6��>)�^�)c�jj��']���=����0
Ȉ�6yS�^���I��'�Q�4�<<d���ܩ��t�K��Y/����vH���ֶ��������
�7�ω`3|��wl��e�Ĝf�s5y_��c�������
���q�s�`4�u�������$Rp����՟�Wk�>�m�k�[�M#�k����B� �Z}���]im�0�נ���i��<&��|���F���w�`d���'|��>|'�rb� [����GI�3ʹ + l�G,��4�T|�c�ӫs{�����1f�Z*p�)e���/p�6�Mw�VJ�%���W��v�ˣ����F�w����,�ƃ�~�ɠ��d(�g���6�&�lj_����(/��N�*�<���dXM=��%��V���~ʀX���7.�
xNIȶ��sd���^a�J��3��-'3X�[�C��}�z0����Wߌ�G�z8�5����6���O)��ŕU��#@�q5u�!�Zj�D+�at�\{�2t�	 �Ѕ��/Y�4�#���CN�V���=5U�܎x1�eU���0�*��M��mF>L�@�q3�K?�`�3�l�c2�����^�@ӣR-����5TS�|�_�
+XR���@��R�S�g�A�p#�+W
4���yo��/���G{*Pԗ8�Ó�@� ��+H z���-��ϩt����,�LB��64q������N�����ӡқ�כX��xU�e��	��)qۀw��=�*g�n���{9��R4bB�H�9�@��ç�e�\�x�����n�ժ��� ={��斐N��[�hG���e�X �)KZ�*��0^����eAԿܒ�0#�-Fj��v<�e���"͈:K�-,��ҁ)'�ə�>�_��纈Z�+@WΆ�����X6^5�qfB�U�÷(�jY�2�*|a���+�<��=@*/�%�)�xVW\3�1!_O�'[zO'.�֊_�(B���L���v�g���ݥ����G��{�t��%M{������[���T����I[�-[����Y������nv3t�����ߍt�R�\���Gx6nظ��[B��L�]����ڷ��\@���z�����#�z�����VF�P.1b��<��V�S�X`����5ޮ����P%yp%Y}V�V�f�|�̹���\t���f���Z���P��6��hb1�����x�G$l��R?I�fA֓`@YR�@?P<�ұ�6�- *x������rxݸ�����U�D�v"�Q��Ⱦ؟=��ҽJ�L�$/�qW����Y
�yW�Y?�Ŧ�C�̑���-_B�G����9������f�V��s�Q�� س4�!@6��xd�+�N9��p�A	8�=��Y���j��t�Ii�]�z^����L$[�*ߴ��,}.#i��>𕧛�7�Ҥ���N�=Mִ�ۼVݴoU\H��/�X;�ϩ��O̗F/��F��zӵZ��� �豽�H��Npf���3���K����|LS����F��R%�*O�E�g��7U�5<;��`�^��x	|qi��V������h������5�7S�G8/*���/4��@�j[(�����~����aݙ���E&Z��,�4	~h�e��o<)�".�w�Z�x�}",�^&=��**�:��x�DX$*�e�B�q1U��r�z�J��c=��dwV��+e�JQ�����Q���B�ָ��{��i�@x{���<W����ǵ�y[��k�e@V�1|~Vi"T{�l&�aճI�5��#�`nG�z�����(���ڰ�,@�^5�T(7%�:�P1;�E�0wl���C�h�mk"�|��Vw�˗��=i�9�D��uQ�o}e대G�ʓ���,�%|k���4 ���H�om��_>�����,��]g��`g�w�fW�E�� E}��ӝ��A0eũ��w�
�&^HWoN�IW^
��D�c�C��H�����Rc�pO�y�ӔC��k�ص��@^Ǫ����Ա'aG��	�OKN�pE���	�ɐ?�2��7�q�