XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��A������O�����D���f��w��.�x����4��5D���-����'��}�����%B���֔�l�c�ͼm��hho�㗗�'�}Ml�|�j�?I=R�9 �|L��s;� ujLs���76���R���ż��~*��%6��O2g�=(2}�6�k���W�)ҋ�A2���=�=o�QV���%��k�ɭg������Ƚ蹒]T�D8������	h�8�@u(�1Y�{��{��k�
w�4k.gZ�?;��rZ�_�F�N̙	��Te���f����X� }Ga�?��=��,�Ϭ4T�76�)х�K�"7��#�I��ތ�n�f���5��_Q���@o����]�F��B����AJ�|����~k��c`�v�B=�9�����:���j?5ō�	�� )��>�O/>��^�UW��b�e)�.�[>�.��%�w�NCВt`���Z ~+R�M��`�{bĻߣ��H�,����OA^�z�G��
��`�����qAw�2ǆ�g([�M�b7��`��)�/���;�(��|�&-��A��JJ�E��#&�߫����#P�
8G�S������6tp��1�NG��D����o$���P�����7�{�������J�kO+���Õ���z�Z_O(GnH;qk�5s�g�xk�*�x[O<9�RU���ҽL�W� �bY^���	K�yri�W�E�����E�y2
8��	C8nO��������(NQ*�]qy��k�,ہX��>z3 ���XlxVHYEB    2bba     bb0�Y1����q�x!�z�*Fl���Ү؁�h�E�����V|M(�%$����݁ ѻ��!+��j���^ו=qD����G��DH�EiKȟ
�u�ɼ����XX�l���m���)	�d�a��;��
ԓ�Q��.l!S��/�<e�-���t����9�ת����ea9۞>l$\���,>?�]XD<��pƁ�8�h&�F��}�:���t��_ʅ$;�N�m'~#��M�D��E,����Ш��Ӆ�~��
�����x��C���w,����w�o���
��6[g:���.���:�Cޜḅ���4I�D\`�,����1�2�k��U���ț���D��U� m���No ��q�	�(�1��f4��>)��mY/���ޭpZ8ߊ�!tG˄�L)d��9ǆa���+�m�Tt�^p�,C��ɢ�Sr�y���� �WG~c��2��74�UKxgY�O��%�3׳�y�cA�+L����j2l�/Fz�m.�dC�>Ό6�vjl���݈s�TQQtO}2��/�n�U��G�E6Q����E](�B|}e&��Nc��wˁ�L~�U'r�sb��.�E��E̎���@?O#���3���(�ǈ�ϗL_�����8�fBXq]���Qp�a�)��2^���ض����	�[�����Y�	;.6,0�$l˖�j���Y��k�P�S6�H��-��~���Y��i��[ME�j�l�[�b�k�	^й�xBME��SZG3��{z&>����Q���Fj*v��Iļ1�Lh���Mɔb�S$%�L���X���K4,��IW�\����]NO
���!���&���O�d�� .��E	�5���ŋ7ƣ�0�����_�I��~�+X���_��ǘV*5=a8���H�SP5h]��Mǟ��+�Q&eL���o#��(Ws�2i5-��##8�h�\O���.�e��FM�.$���uK�Bp�d����� �yX�3�A���������6��ޢ	.Au)Y"(����
9��qrt6���(8p$��_���# ��p%�ypE��5���1����l��~55-x8�v�颎����6|,\����b�1e�q�
#�{f�����䥔�%Qh)ך��s�WNP"}YaQ�}i	m��D�<��=�A.4;�a\����1D�z���	�_z	�[�a�[�7 �3�Tn�d�,ğ��ߦ�7�a�� $U���c]:a�SZ�w�T�Da.ʥyi�ѳ�d����c-��Ȭ��MD*��)p��f��,�݇�R ��*�I�����,�m�oDzV��k6r�>��?��~?�O���;�c�R�l�&Pd�@f�8�1�w��֊��|u(�l�
�Ue�_�Z,�V�#�t%�_o�L�J5�3mr�-����v��UY ��zNb������a�e��1;� *��.�f��+�J���zs{ZrR�lӇS{~[��J�F��f���d1�{d�����g��0�?���Fl�Y��K�+z2������C����>��F��&r9ј�3A �b��v���4D��ՈP[x��9$8�8MSp�}g�}!\*���Cr��Z�/�T�^�at��~	��tgS�<�I���o=%ƣۥ�,;랂�X.��~V��O����ʊK/��X%����%�h�fBb�G�������8м���w��y-tS>���;&=J�Y�O.y*����tc��.����^��.F󤿊]�(eR?k� � �� &�К#s��]ʎ0h�8ͻ���rw�*���M���m�$ș�|��XOT�J���k$B��q ��lg����k�߸����V�D�k�@f/(��jH�s��˷��-h��{��5�����\n�heB=�_��F��c܊w˃��q�Eao?��,�iZ|��*��M'V���ɡ*�Hu�FmV�52�XY5f����n�}_	wf �_T����8Z%��_��hWwI1�>���{cPt��2�#��D��{@�'c�]�ή<Eг{�� mnl��6������թz��Y�Re�-�ze$z�t�A��T��U�N�84�x�س��N]���m1U�v|�,�<w��M��=����vV+���sGS�F?Oq3��t-E�h�����K�PN�ʌ�hy�Z�9���d<�m�/�h	%��@�;:��U��Z����0��)�2��M����t�Ǒ҃޵�iV�{��i�G#�5ٗ��l��0I�*i�}�����ce-��]�%
��Gq� @�����s��9��#C�g-�Ԕ��7�M����੡���!ܢ����Z:81p�U�/�)ѐ����:6�s�����:��n�y� �}�;c��/	Ӵ8�ܘ��L�F@���D`�ّ)��=A��!8k� �R���=h!Ӻ�bm����a$e.

-�������¨���:�Ӹ�V�6�+#x�W4�� �� Q�&��p ���âڶ�IR�#u*�㴆[������&"������C�� ꃶ��w�p�Eq�A�"KŽJ�����5(OI�(c�wr��7�a�����^��J��hw�d�#(/��I7 ��Y�������K�fͯ��3�0G5�!q)�ަN�~����X���֑؏(��s���X�<���c��HҨ1YA�E���p�OVL�[u�[�|�,�k.ǁ����1�F�f,�`(��Z�]�W�i�a�t;{�gv�.�q��X��=�յ2;����x��^�k �@����mn{FD���_�,�1o]k���u��s/�Cߋ[[^���X�T���ǒZW����,�c膼���x,N�������u�_�"��y�翪]@���>4��h�N%��U�V���"��l���8��Cf�Y�Y��n���i�G�6�9EQ��_��E_w�������y��T���ח��Z1 x���.�J[�kїV,