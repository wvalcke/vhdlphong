XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���2	Ĝ�d<VS��&����5B߄D�w�zI�[���tQ==�.��^�l{W���2A�.U$�h7�8���x�_b�EX`�46U7����r7��xOk��k��VO߮�ƥ��ٚ���ȳ��%���	g�,�6�zmI���ДF5�~���i�U�C�;��3���T:��o�XF���N�	?��.S��/��
 Ye���	�k��n+�b:h��Y�� Tͮ=�{>.@� ʰZ�`�1���'[Є���8�,Am��9�7�c� ��E1Z!��p����\���V3�����tm�����GOvҷH b58��ջd�'�}c����"�s��i�R�4(��{�����Ҵ$��g��Ǉ4d&���bc;u��ҟ!�	g���Q�!����ZTjyd���d!F ���ݩƤH*n짍y=W��6Ц�7��@�A<�C��v�CTJ�6�����R=0����hb\t�4�a�y�N�S�T����V����}{��&�2��CĚ"�i�z�s�F��
�A�vTPE�(���L�͸/g:�w����>�?ŷ@���I~nu�H^�"E����X3�bQ�!�#۰�a��%�㖼�0h��.!���<�2O�_�S5h�͝�3��l�aDg�Ko�TL�g�p�p)��l���D��N������8ū+���1���cֿ�~��G?���R��Q��0+�U`8i0fH��!�Kxnr�b�'����O�ڈK[ʕ������$XlxVHYEB    5e75    1150De��VFO	l.�׋:E &�M������f��Bm�B���
�v�
��*ݶ�+���佣Ġ_9�Ḧ́\/�Z��W�?3w���w�Qل��;�awe�ٔ	ص�6�C&j<���i�����."�6C1�7J�HG� �bM���H��u+9�ն�oB�B�d�$R-冬Q��	�k1Ys�w�g��B(<�s��U��؉�y��cnY"�0�%5y�͂�+�=���?�z��v�<�V�)���2��\�s�u��U�Ҩh�K���u�.B���� �#:5��Y��92ys��\�S��̒�5`vn��f����u&l�VL�2�{��2����C���R@��V#�NX|;��?H�=���|�,�K�sf����̗�uZ-�_���{0�f:�u����H>i�/F�"����K`��-��mxh$Y�
���8đ�(9�m��mo��zW�E����}t �Г� ch3;m`J�9d&z������Q`٬g=׶�t?�-�# 	&G|��}��B��D�1T;��,Q�y]��S�B�O6�,[�%ب��sL��w�J�z�����jc>�3pg�~y�����O�\w��5%���S�w������rŦ�ћ9�ش̣�]<Yq���=^/�F�c�(2<?hS�  sѠ�z��mc�x�Q׷��!���3��K�%�1N�'`�� 0�c��a��D*�o��4�j�����Y�&�����Y��[C�t�d	v*~��s�=�L���L�w]|,"8T�ϛ�U~������%w���}-�q�6��9�!?�C���#/��N���x����@�,7���()�(�V�$XS�^��R�㟏T4�m~u��,���Vz�0�	����%@���𙰏���/&)��.ד@N�b �b�l���TKu|z�q�PS��*CĳjTiF�+���P����7�����3ڬ��<����T]e��NJ����W�L&���,z̬�8�m;;^h%>j�� ��Cvg�v��D�^�L-�s��&A�VaEB��x��xV�9�ȕ��9�re�暈�3T&�G�B9�v�����3�p:/t�����W|�r
y�%[��삵p�e6[Q�"�B�n��7�Bc'u�I3!��"E�R��!����n8E���-��X�Q��{�����q�c��1�R�UX��f�/p�� ���Q��=)��ڪ���ÿ�f��U�Pp�޵=�(���-=t\Nz���C��:�Y���U^JB�P�i��Ԁ ����9p��f��(H��eV�����L�{%����c'�
���~ĪV�ϥ�	<���&��$P�ɼ�/�b�\������@�F��ܧ�n=���?T�x�O��ᦜ����c�P���QgcKLD�����s�Y�pzxH&�A��M�&�h�	nA_x�0�Ct�����\��[Z'��$�p�8E ���αq�]%:<�_=�����hvV"Ůa>*e���C�7��"n7�kn���߃��?':b���
���]U�Y 2N*`DPؒ�����9r$��_G��X�uh�K�ݴkr�i��&n ���n��p��V���7S���m�dfQ�Z����m-@�����C_����q��]��#��T!/�g���3�`(�����X�=�9.�6���#�+��~�]��7<W/hQ�͚��'sr_v4d�6!��H�r���
P�9G��م��(�T~!ė���8�3
����_w�=:ܴ1h�?I/v#��V)���#1�b�n��Z�a݆ױ���*P��/��W��oꭊ/�/�/��G��zK3{��VZYF�}�,���4?�6f4�qø�v��.��L==��.�6#Eg7�I��j�"�#�I�h�j��/�_	d��͎X��۩��Rj�my��%y���F�u*�.rt����VY��ˉ��1���B~tl&5AsI�T�	�;���" �0m]FK0QG�'ONl�<�����N~r���J�/�V=�n��FW="ij:niQ�͞��8Ҽ���2C �\�������c����"YV�bz�#��*v5�4��
���Q(��	�褚�j��{�Wfe������k�2��{B����k��#�/�儹�:Ob�jµ;zMd�Ŧ����T��E*X��4�G�Y�ߍĴhc`e��Vb�s�y���ڤ��6T��Tބ��,�B���4"�����mH�a��`����F�]�ES�)/ą�
0B�����3ܷ_i#C�DB��,��Os��x�j�FÐ���ح�I��H4�}��"� d�׵ߦ����=��(�\9������cd?�3=\V�F��s��&>70$��0��m��TP��OX��KℯQ��kb�Z���qb;�ܗ�Yo����x��e��R�����8���������k�szI rJdA$Y0}Ѫ�~���fq�/RsL�NG��!'�
��N�;��V} r 9�ŧ*���s�ٰ_G50��9.?b>JB"�v����m�~M��N�Y��-!I���Y��!DQ�L#�kh�
f�nr�[h���m���^�}	�Cd��q�h ������|��#u��@�B�]G�~۳��o��g�k����� ����Si�R���İh��;YGk��VSox�&����h��m� A�9F[��e�ُ^
�a:y��@�!C��(W%�eJaf@��L�&�1�u�͛�`X$Xx��!5�Iq��*�G>O����%��}/�Ǜ>��*���JU�6}h]�]&1�H���7�@�oV���n�x�y�Ҟ�lq��C����Sa�N-����KPF�'���1�0�=�TJU?��ō��N5��`
Γ&��N���̚5���W��Uu�Ήn֤,'m��ñ�w�����fϑ	L	���YB��`]_:�Qk�q!��9"{5>��67'OZl9D4�	����g˯����VU_}�xh��c_ߛ^1S�gԺ�� �w�#yF�kz!)_���.(�ھ�|�%�h�ֿ^Q��Ʈ�Z8õ�<]�7P[-��g+j��1�Ӑ���[������q%[;��hࠖ�q��jk ت������uwE����v���jt�+�A��~b�g,)�jԉ�����c�u�e�
�	��Rw�������? $��0����L0�׬R�j�!6���}dB�A�e6J���b��P��p�S������wi�D��'TO�4[�i0�C~j�'yБX� YM�9_�y���hc�lt�'�����4��[�!q<�s֭;SI��n���t�5��_`���Wg9"���L�@�/+V4�\��j�i_�Ղ<��+�;)U�K��֟�:�o�}�2�+q�[�����H�goPX��ݧ����=��m���+�de�}�r���s�o�Ѹ>����M���J{�]j�Y��2j��n1� Ec	��6ᒌ.'Û|b&��c���U�Y�-��t�N���Q��6��;����˒^�|b�z6����Bi�2.Q�r=Ý��� 7��>/��#�$�3|�u=? d͚f�Llp��]�I=�[����Pjf��@�i6iL��/%���_��8��-֢��m@8�Ň�
q홢���S�9�s[�Y�$kp�7�����BH{񒛾[B��]�*[��;n��d?���06�����in�<gS��KVT��Թ�_L6�fxE�)�M��+/s�L�6�Ӿ��U�����v���M|C��j���p� I@V�1;�j
=o��̼�|�] *`k����ƛ3�C�U?��i��O�YcP~Y�O	����2 �
�aw�n/ب��J4��(C���o��ݛ���]�\g�J<e8�!�����n�Zp~�ɬ�(?N���5�7+�A�@ϳJ�]�#e7:*�\�a�;��?Qk�mM
 ��@:�	�Ѹ%ma�E5���U���`n����iP���mj�,O�'ٓ0t��0�W�dar#x�D�5��� we<���D3Q�ph:�t>B�`f�'���NR)�<�O�����޲�y'\��V`�x����PS���%Q-K�+�z�������BЅxvH?z��<8�'$��f0G���V2�5�5o��"�8����B�~�dnE�������ۚ3��a��nHv�)���8&��2���ǟ0q��#�ٶ߻����BM��E�Z'T�>v�����51���T��ۣu�qO�z��U#3QM��	Z# �]�y��*A8�\x���4�ӂ�}!+�R�&�>^�VJ�+rF��R��Ebm֤�t>��*�6&=}a���E�<ؗ�>ϖo�PYgxc`����4�;#������X�I�e�~�'�