XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Dð�b�����	���fAvC��a~H���n��Y�Y�Ekm6��
�j=���̲��l����q�*�h�\?݊����T�v���+�$�3�=�2)3�GI�{6�M ��ܨ��i�/'��������2�s@a����qZPNA�H�D�j�#�j92���~260��)�Z�U=�x#�ڳ��Ѫ�v����k,~�~���]�i��&0��8���x�8��X � ����<��r�g?K�LY��	)7���h����"�E	�.!l/�6A��X )�b���e���n`�()���Q-"��eOj��"%�Y�;A��6<1�JBn#���,�wmd+�+��E��ō��%[�����;�oSF� ��	��Ķ��.��KB�Zm�,ڒe�dk�s���&l`��S1%<~-��:���ʉ�*���9o�����(����D/���頬B4ʑ�.���)��驡�n�y �a������[���Ҥ���;�G�ƽ/�v��E�����,qǥsz]m�R;@M��
`��v,�_�(T�6Z�9�niW�S��-Z�C?u`�P������[�R�bs/�E6&֢6�-дlI��>P#�W��rk�N~U��I�DE���v+��O��ai�W���:�A �Ң�shF��1��s��|�����KG��E�e�K��)-m�,T�|u;#�ʸ�v�l�[������,�4����
I�$�T/�$�ʷ�`�����YR�+�����t���`�Ih�=��XlxVHYEB    2bba     bb0]znt��\���a�~�-�O��՝>�!Gxp���v+�䧑Lb�n$m$>r��r]S���P���-�T�{o�Lz@(��ǲ���60�^d!�����F��je5�k��>7�[5or^7���6E�μLSRѽ�9��8����JF��j�s�n�_����F������*AS��s�m���GO�#�ꅴھ���Xz�}���B�F]�3��V���p����2gL�n��2Yqb�e�� �[�G�9�JO��"�Ƞ5M-�T�� z�qp���B`���l�3��Ɲ��ѿ0o::Z^�)���~����3�0@$����Y�b&v�4��i�L�Nƿз?O!���"%Z���]�w6��CB6���.l�g7���t����Q]1v{hF8nHk�}?��ʵk�x�x}GMt�n���D�T��~@�5�w'2O� Czj��+�]>����Xz��q�,��^�ʧ+X��B�����%� dVZEQ�@���E�Y�G��FY�?��ʫ�L��`�� 럆>
 ͬ���n\�L҂c��ez[���ܼ����O��p���k��	��2뤬�|�M{B���-Ɛ�:6M�q�-R��Vt�;=K�	VO}T���������^a���
�[Z/�*J�y.ˀ�����8���
��,��A�q=ʧm(��A���wE�O?BO+ϫ��0^�f��>�K��Rz���4�ʲ4 ئ6m��/rf�S�:��<����HH�k�@DD�)��_�pt�3?R*b�t�Jr1=/{��N�Tf$��(�\�C���(�I�ьٌ�ð@�0l.��6�Bz SY@�o���{'b�^�u�I�/�]?�����[��_U� ���h¿�G�W)�AF�U��g$��aBh��KP!���[r�WѨ��k���šn��~9w/�4�#�P�VT�oa�"MKj�`Iʥ�I�:�ex��^������͔"�i,DA�AF�5�D�c�����ů6�fr�K���Q[��͛��ٚ�V*�Vr\B$Z;�l�T�{�
��[�l�8.����Ŧ&>��Q�_���@~>q��{��L�'<|9J��Rx�P���Q�r9�!N�w�}���m-���2�)�ee�N���\�ʄM��w�Q�a&.NY脉[f�A�#G#�>e=��p�ݛQeAI����F	�w�j.̸�{����k"
e\Z-���e���}@��&3��_�=|���=�����(@Z�`����쳂�����x����Њ!S��8�C����`#'@�w/��L*�OI�
���يЗ's���1�����hNa��q�Xk,�����}��(Ö��2oG�]�`��IȦ�iĈ�� �����z�~7�������ģ��X5�O��Bq�meY!#4��Sq��M��
�Vc�t,�h_�{�v�N�x�����]?�O.�!��䝒�F�'T_B{�Z�dP�u�~&�(�<<#h-�>{���4
�&,��Ljk>'�H�	H������T3�[�h]��LT�2y�3՜oWP(�Ed��S�E���͕�����������K�!
U�R}T0�{���Ai��ƕ� :��C��Y�g�#��4F#�$�M2� ������(6�X|�6����:��ș���	j���s?��t��:<��v[G�ДD^ �]�<޸xl�,ąj��j���aI�{�$�D��ze�����(6�/���D��ځBAAL|��$�&�
�m3�mr������[P
��K�2���f~�/O��?ȃۭ�.m��'�Yp��2���V���'�n�S��lI�rê�Y(����l鶹���>�18ީ�~���E=�-8Q7~ؗk��J�#Gdj�i[:�k;���
P�KEY��?6���h�>t���=�(!%����;�k�T�����O4�cTG����d�)����9/L�i�~6�&hm��E7����.�숮rW,��=`��n��7��w��)�w�U��)q*�˒;�EA=9fBQ݈��]�5���Mͪ�#Q0W{�7/�ӢE��,������y:�������kb�R�r���:ڝ���<"�O�a/T�t����T�	����P�l�U���������bD�=���3zxU�3���]���ED�%�bE��f=R䆯phy��X�b�6�4Pb��ê���������%ǷE�Q6�k���:O��&$�#;#{*L@ǫ򧷼Z����t5p5���uo8>�B�hk�W���������~��^�ڄK��T�Q����Y��RN�7l"�Y_}�:4.�y���W��~R��-\*��9,��+���c�Щ�h�9�i�sKawyW��;X8���K��9���S�gY���R���.��zUY�M�=�?�k�K��I*�:	x�$�����D)<H&9=��S��<�l괒=�_W[J���1[�AOTn�%�Q v2_�Tn�6[�N��|j�M;��֧���@�����������1�7뗴��`'5\)���>�xTg�w㳳�.k��� Yx?Z�/�<�g�>Z���R�(��v�DN�F"�jM��⃕���X���)�Q���LT}(�W��|i5��
&6j*�@t�puP4%K���{,v�#	3]�m�ڻ�ڶ���"��<H����b���u�j����HD�D�k]�].F���b�K�����[_���6S��wZL�͘�k_0J���zĔ���g�䍐s�9h�@2�-6��\�ED��I߭],�U�}*���w��4��z^nAi\�d�Y"��+C�7U���|}����/7(xU�0�t�k��F�@N�p ���kerJ=+xZp�cA�K��S��TV�w�a]�C�i[U$ z��xw��S�� @�w�h��
�M��e���C�51�IO~U0�Ux��ÄKO