XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��9;�P=���n�1�r��6��c�C,��)*�rGU�ǹidP�*�q"�e�h��Է�f7�N�hB!�a�^��l�D"n�L��uv��X�i���poH�|2���vDv��6���d��z����c��d��po�����G�j �~d*���X�B�{i�)�#�f����!�*}���zG��R�l��+�RL\p� x�+!�hRS�1v�d����rb�����Og?�Qמ&����'�;�̍��IF#j+[֨6d�����|�|6��؆7Pv�bV	����O�+��������{ذ�t��@�]#�,/��K�f��m�U��Jd^��U��p��ӏ�j�pb	[�!��N�k�?������X�J(�}=ˀ
b
�}�M�;�B}�s3Vo���Ӥ�%ĥ�B�<{�k�y��(.95O�l����u���R��4�~*���ƫ�"��Ju��<R�pu�͈��N�����/�f�w��lj�WU�/���n�1��h�@Y�]SOz�0k��V��i߇�ods+<���&�*���{l[`�J�1���k�Qs�_�����&i��)�V���5`kGFS�q+$���* 8C����R�ϹН��{	�	�)��4������a,l9�lйB�R�p���xd��ܪy��ҭ��C�7DZ���O%`��j���_ҀIr�#��1��ٲN�B=�(3i����":�3%�zQ��)��*�r��$֡�ԭ��R�'-�4XlxVHYEB    4013    1050	��]�h:I�����4�A�Q�+�]�/�
�b>s�O�2�g:���c�	˺�k�>���
:�sR����p�=*����5�z�qj�� _g�a4	�wu{`k��cc/��
a̕p�#���/԰1�s�3����R?U�xٲb�����X�K�����@U:ꗫ�kV��O�*#ԈP)J*��K��8h�U��(��k>�������_�����`�=W�L�y���,��PL���6�)�!	<�C�����E/���_�'B[��S��� �O�/��!߶����r[���H��&a���_�����v�h�i�A�u-�\x+MsR����od=� 7�,肦Lz�VP ������iƼ�#�#���ܒ!���{$��D��
�;)nT}'��x��O��E�������kL�f�Ar�8	f���4ҏ6}����/�AM0�؁Vo.�
�i^��Y�:���"}*��ʳ�[�<n)Q2�g�zԶ�1Ț��v!;�y�Rrt�|~��"4<�(�y���Ǵ�.%yEޯ����P�[�ܥ0�.�u�i�Ña���ӽ
&<�3�����W�����D?���
@�4�78Uz	�����܏Ժe��:%�e�w��
$׍LM9��2z[�%ɂ�+�Z�tI#�m��G=oUx���t+Ch����_a�X6���� 䓙p����"��.���=-{�_{� ����LNR�!��, �Ժ��[!���_��ʅL���vf��M�;�^κ�zx���(��$k�'-���n��J��Ò�SN�-:z�"P䴐(���^y|�V��5д�������Z_P�V�$_f�m��U���^���dڈ�^����,w���f����AmI��
s��@�����d�P��@N�m��D)���#ݡTl�� !\��@�$���;<�Ļx}I�夞�?�e�!עZ-�^[�&�h��@�?��=D�u��	5������,��G"�����/z���[U�Z.\�ٶ��8Q��c����:�6�@��Nmv؈�A0x�a_,���:o狥��]�����i0�WHh�VP�-�`�̅by��07��m�W�S���%�Q������㗁	�󌶹�p��M��8�����3cN�p=�-R���{�4&X�Q86v��V�a�g|��W;7��>0&��%�Ա�����V�>�����塉���t1)C�i���	6��h�����>od�[r��W���	�Dж�l��S�z��z	�m�Ǹ8�(�!��Ƀ���j(6�z��1�n� �&t|3a���
p�4�����z8E���w�5k��z�o�ŷL����H˂��8z�����(��i�*` �,���F׻��gf�%)!ΑR8���.���Q����[��br�'I��J2����pq��$�'�g����Tz�qt0�eHy�x���&�rTx��Ը'T������G�#Yr"�-���1��bid�Z5�
����z`MD8hd%�*�9�=Qn:9x����Jd;��<'��Vc���aV���Z+$��w��3�tؘ��S�M��l�j	�R��ʙ���E�|�\/�(�Ō\	��Z����o���d��l_��H���yO�w���uc�}@�8��X�w�|ti��n���3GhɔT���|=�`5�O/�df�y4KlvVP��Y�;@�ix��nK*��x�C����7�y3wjx��Ńԥ��v�I��I;'���>���]�>+azZ=l����G��. �dq/dBo�=E�"-V���N_��a4&I���T7r�вW�^֞���Eu�-�~̾ ^�J:�uŰ�����.+��3yŏmj��{-C�C�G�i�97Ұ!�c�~>�|/�o���>,�n|����ъZ/PX��Y�ke����cN�W6O�9�p;Z�8\➰�fp��H�`Q������T؁��恇u�CBщ���E���N���~OZ	_�VP����q{C�{u�ƿ[��L�d�=k���-`6u���j���%+����QQ�\&[.3i3F�'�p�m�!h��ڞپ�	�&)'�yLՇ��)y�@G���"m�m�=���6U��De�0��2JbS-��s�O�؀L�<�@�?�-r߫������QL��q��+=;@rU��~(���L����k@�k8	 bb׶s8��!�e�r�<^�_>�w�]���h]��c�b[h�	��r�!ޯH����Q���YF�h����V5�H���\���#s���Yd�k>�[-�7���eFK���S�j�Џ���<�����4� �����%k��Df_z�{�<������+�l��	�k迴�o˥,t_N��[�u��*e��$�Rw����]�%�Er����{"��(�'~����8�,��t�n7櫍���N��t�֎n��@����׳*Q� � 1�5(\iP�Ebaz�h��\�W��X2/��8	�{����>��B�NN�n�2qn������e&��_�]a�����JDi�4��JY�Ŷ���d^�C�(ch���q�+��eP�:J����C���MF�b�c�rX���[b�A^V�..ʍ;[(�$�U��)b��fI�W�.
�ܟn�~\o:Vw�w�S�C?8�4y)[�xyU0B���h{w���N��(ɠ�h�)�	��8�����X؄�e�� ӝȇ�x�0�r@c��5Ś�z�[�O��}r��n��vrԈM�T*���YW ��{�+���zΘS��@�LG^���3���;�F�8�S�a�$|��H��w��Y �Y�R;Lυf�˘�O�1F�4#����p I��G]r�C(����N�J�s���v������x߫������硑�PXHŰG7&�PɌ��n<W˂� ��P��Ԅ���$5��Uc�g��d7q��:� =yUʑ���M�|�(H��8_{����T&���>�����ԙS��R�ON�s���J��>J� �{����(9B�_����P �8�A�n%��V�x2#��g�OGL'��Ia`:����5���7 +�fZ���/p:��35�E{xI��0�́`D[�bg����gW �|.�9���,\g��-�f�����K+�'�~�.���ҚT#p������J2s��`ݳ�<��%��QJ�<���,y�l�iO�rv�	���0LBRp:~�W�>�L戞ѹ��20ToS�A@297���tCeu��<�ۘ��_8����\~�[9�ǐk�q�.��b�#�<�KX���x���JJ�#�a�X��4�oͅs;��^pL�υU�)�S�!5� g'6!�@���� ;��^9���/�b�Ϛ�������k�"<�.�~���n��ۧ��+$K�O[@��������ć�:a��wb�!qN�u˟c�=M�=s���])}��4e��Sy	d�:�2tȘ�+�W�� +����އ\�w#%}n.�#�X��VM|�æ�@�f�
�VJz���Kp{��|���Ù5��=CtF����
�B�w�Q��M��賲�\����%l}A��3�)�.��L*���)��k7�('S���+�Ȑ�}���7���,�/�/Lq/ز�T�����vVdn�Yo������H�~fpđ��������ƪ��I+W�]Ƈܛ��FZ�3�-M��utz���a~;��8�po%�k�����H�SeYL���1�U�f�D+hga0�{*n*���R����(�e����~3)R��4�+�b�~�>��O-¨ц�~�߯XWֺ���~����h��`�+�xm���T�I7����Q�i����ߍ*���` rO���A�a�t��NB��
�.�!y?�{��z��~�n64��U���'[���6 �d��8㩶:�t�M�����:܉E(%��oo�\YwF]MI�4�}8Ru�FF�U/+z�7�ѴO��jVR�����z0ܣ�x���M �<��G��g�]P�=%e��)��;fY��y?�%v���L��7? +?F���Y�)ν�I���