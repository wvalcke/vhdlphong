XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��3A.`c�Z�5k��*�-a��';HL��mmO��NYN��ؤ�b�'��qv'�m�$�����=܊|����ű���x� �rn���33��Nj�zZ�{��Q�ۊ��
���.�l��<�{dm�4!�\��J$:�_#P�i=�W�Ɇ��:۵ XZ	oҴ� a����	�U S��ciL��%K��]H,�c��Bo$�.0�����+���(�k�`�)��"�[R1�M�ý��/A����[줫�?_��+�h���x���!ZY(a��������/��y�ᤎ�/�N�@�%ZQ?Y9���w7;.N����U'�7�sE�=R�;g���_��;_J�Ɔ���bj	��3��1��g@�W�/�8�����4ONΪ)�MŎҩ�/@xE�nbm��;@.Hv88�o��br���E<0������p�ie)ZB�˿M{{��+�4m1�XCw��Z�"������
��=��߀dwҍ1�.-�c 7W � ��$���\վV�TU]�S����ͭ��O��21�F4�.�G�ezVMIH��T1O�$��`-��g�#����+$;=N�(�����.�j��ot��p}Äv�������?�yH���m��42ӰxY�de���G0����Ȯ�i���l��)��>�*V�T?= n����=]A٠�@�W�9V����7�qޑn�L���������W��{�� `�������mlŃ kQ��X6��X����*m��|!XlxVHYEB    4ba0    1230�Bң���,�2Ѽ��r��F������x+�q�m_<��YY3֌��R��o/�-�0̆�����G�����n��n����/��2�����1:�V�c�$��e�Y&�YĀz���D��'UI4��B��qA��T�\�jP��FѺ��0�&q��?�O=���O?^x�`��j�������}����O��8���X�H!T~OS]<6�'�=���;eº��I����u���l��fw~�xY�C��
��m���H34���*M`�
on�5��n�[:��dT�>:r����� �Z�$�c��<�]`��j��#�/Hvz���B-f�z���0"4�r�d�3D/�%���w ���
����j7����!�K��PԴ�i��J���k\�����6�N��Ř �,Ae�~P}%j�k�C.����>���k(��k�c%�Spjg)�D/��,_�2x��rY��qM��D��圠)g��M;�ۢ���#��X�%�H���� ���`�����ӻc>�:����o[/�m�{a�9hY�w�#��wŻ�����f�'�ɏTӬ��,��{���W����x	�]տ�o:4|2X�VX~�Xo�:k�M��_zO��a�[_p��q�H�5��Q"�q5k6V;��������R�n1�¼4+xp!��牎����ϳ�zˆiS�}0+�b	�e�[L}�����A�oӦ��d��oaN�۽����Ow��ߟ�D�E�����ўu��h,U�ߛ�v	E4�4'f�bp�(��yyv)z�'�0��?A(�h�50��	]���ܤ�̛�N��	�<�Uzz��h-�y��1���)���B̼�ߠ�^<}X\�Vx�{���1~������L��Bv�����?|J�o���}k�AWX6����e�ِ�[x�'��RP��.	������"�0<�?����K���a��@��3m�!�S��I���1l3�ۅw�͙r&����[/o� &��VP������<*3�W����%�һO��)68i:!��ź����$�辅%b8�;�>�����ܩ�-�����QO2��
�<oH�-���~��]��ƻ8�"��A �?��V.��vil\�ő��|vL2p4�>9����31h�3�$�D�t��l��/0�	�<�&�m��d��΋�W1�.�Hj*O��n,ѓ�v ����@��� �e%ݽ���apTA|�Ge�.�M1� ̣T���d��g׽��TLa�j���'b�.��\7~#v��S��@�����{���%���n]�B�����1A�G�f2.��%r�������We���,4�2���@h�-�4F�<���'>�����k����n����	���E�m
��ݵֽ3��zpl�~aIB���EVق�?K°>���@�¨p5ϋ��4��v[�&O�c����HP�8���r��s i>\��Է4�G+���b$������\�����~'Q�+�S��$q��y�25��T
�<�L-ӝ%?�}O�͇�ú����,{�f�p��������೥��������L<���ʯ/;���~=���Д�̤N�R��`��D͆��q��/��x�)oRTC$����~���Y�>櫽����HJ��¸�[����:MK¯�Q���/0��y�PPx���a���18Hu�v�p]�Y���9�ve+.��BcY��9��h��+���5b�E�8����Fу�67�?��!�.������? /ؗNɧ@p���8��(�v���r�o�95��kLU��ߗ�7���7ԥ4�_���n���4*�ر+O0rӃfwDn�ҹ��Q�nV[b�Z��j�ٜ�`��'��4_�L.�pS�U���y�q�<kŸ�zs
3����H%e��e�>̝��V��^Ș��\�d��'k���#��"xU|h�� ��vt1W�@��VT�/6<5��Oqy��Q��̔|e��"��5�G�PQ���o�n�ܡ��U0oEf��?��f��H��&{i�f�Kj�f�qK5���/�8�R�J8	쿡z?����x!�a��{=�U<�����^�����O�gE�q����c��Jb~���$��x�9ʟ�R��.���q�c���*#��8E��ǻ,ǚ�����
b��A���q���S/�Į��/E�k�@�ՠ�}��'@־zr�����2���a��7&�H��vKh\��"�^�O	�;����O���4*���DZ���Λɐ��xv�і�}�JX&��_{G7�|?��>�)�O��?q���|=�ǏDL�Ss�4�L���/��@���&�'��W�Ͷ~�H���22rW�kH�����v 5�-���ed���X�a Bw�*�����w���1mޝ���^lG�מ��TK���`!xѷR<;���O'��r�-�}|1��w�m�q�^�����������RC��,s�3x G����k+<���� �M/�ABE�}1��T�D�1�&�*��۱�QԚ
���&�T��_8�|"�f����%�GtD��}�Y���$����%đ .J��j��3q;���z��/��~O��Y@x���Ў9�^%w��Y�2�O�ZJ~���!C5[�RY���fg#��̈����B�mE{�m�g�6�.2�h�9�U8��\���}
�B�T������ٰʦSe��>Ł���.�qk��ӽ��WZ�܇X�rr�>�NO��r����s �TB����ǥ�v,�'�YcJl>�z��9@/քŉmm>KnG�;@R� %�x ۶J���*���'�6��d��ce�2_o��7��Ex��a�'�i2)U(I~f�EԻ��w ������~~Ȗ4�)�{7�d�Y�)��*�kzf�
�Z9xJ��OF�,�S\yv�d-�ϵ�����3�|ۗ����w�ַ6}b ����H��q���j!��T�� ���Vi�r?��!#�)�kG9�	JyO��:�ܯ~�Lc}R�6^r���l�I���������.2��{�B꒳�i�D0�Npw�Ϝ�V�4��8�b;Sh�@m�r���=(c%7�f���l�ݔw�{���p�3=W�����������p �k�f�bH��N���lDH�&Ok��@�yz�)�j�|{���V@���OD`U��roq㨆x��&��Il�j��5�P3ʻ�4%��-aG ���ϖ�v���U��_��IF�/�_����0/x���������j�>��Y�k%�-����0�8�}��ל�q�Ee��S�纁��5���u���I�/��J�p�O��&��'��T���~������fZ��!"F����I�4)b��7�t�á��q�����r0��ud0P�o��fd�P���ܾ�J?����N�w���z���F���(�� �t���X�n�w��|�j�u!��UU�e]���Tn����@ ���_A��$���ᩋ��1V]��K���!�="$�4�]����h�آa�����$x�6�d�D�e_����|��H#�1zV�P���^XZ,f��)��~~`��%��}��0�L�C�WLQ5��}��N�a�l�ܹ[V����-Nx>9�J��M?o�U���N(w��W��қH��!�_1����_S?1�3D��R�'p+2@b���a�X�ܟ��%$�8m����~�%d�;����<�M�SP�냰���-��f{K��=[�V��M��eJXc@T��6�m���5=D�pSI��B-��
5�=N)�z$4eT��Q�ۤb�%�u�G�'�.]1��:�P�t]���u]����IvRؒ�w=�&*�0cng���<q�!������3�N�OD���}�!�{�(M*������J�d�{��w`딨��K�	oc{���,�M��zľ/��Sy=��K
��>�y�d[ڸ����S'ѿ`u�@ S׭�|㤬Qt!)���bI6����]��'��[������kj��KB:RS����c��@�^��y�Sg���u�k����ky4�ГM�a︼(��AMR-(�S�"��M߭E�d񅯎�@Lmo8�� ����3r{�P����i4�4�}�N���;��QDh���R��d�!�A���FJ[��ԴB�W��t�r��g�^=�xʓ)7���n��:��C\�����G:���}P6�Z�����W���^��'2�ق��D�CF��@�;
#��c�/���OE	��īY@=���|���\ ettD1�c�<����lrCE{��*�����֜�6�ꃬ�Gs�ř�
v�ә쓟 ��໼��!t��	w�8���l�:�������� ���-���i9�a�'��8
���PH
W���CץTЂ,&���jٱ��S�▉���D��(۶~ [������#���K�3C!�ƾo����P��gy�y5�s!=�� ��s����"�P��f���r<�5j��<�����9]�_���]���	q1#o�gA��fR��j���}�V/rȟ�:�m�'A?��Y���