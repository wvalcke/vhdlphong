XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��҉7�$���b*�qF�+pc�k�4����X�؍���I΄k��?�=+�^ƌ�1~zv��y�V�����.�4��BD��9J�n5͊<�
�Fǳv�%��\z$�L����o�0����A*7��D�����v�;N�vց����أNs��9��"��U�p��*g"hq=COJ.��iG����~GtyZ8U�o%U�_��Q�����0�2Rytry|yf�z�,"��J�'�f�L~���@[��;~3�J��tg�AcMʄzl�c1aQmK�ǡ��~	M�����웿A��pՁ���4���d��~G����%���<������8x����+�dvT��*.<0?r��^��
�4L��Zf����[	��Ӏ\�9}#~��-1�B7�P��s���#��l�D�D��,Oorը��ZsʠO�!��9���è)�V&:�$	��	z��"S�#���?�k��r�龚c}W{�k�v�pAמ��70��;�=�zc^Xc*�{�����(�"�����`G�T��z���6Kf>��-���`��Ժ����@&���d��Y4��|3#.������ОS�4�d[��E����C�Ye@����� B�!����	�j~���Pa���m��v��k�8��
����ݰxV�Mq�Z�>�f\��i�X�\D�Ď'�bݣ�>��Bϧ�89tk�U�^/d���.֔�0�̋-���s�����X��ɀ�|ώ3��v�f�.2��!��D��wt}c��XlxVHYEB    3357     c80�X�7y�>�]���+as�RX�p���^���	5
�Z��{%5Ǥ�?��	�p"B@ƽ�����(���<���5qH�y�^�=���C����6[�*&��J���w�'�:��$���~��8�1-[\���4P�O�b���U��W� |]6�gyL��7�m��¿z���.+/=�F�	��Ԃ���ۧvB���1�?<�C>�t��b�	��"��ݨ�+�
���=�i���=q��6����;ܵb��K�IU�N�~U�ˆ��S�^:Y4%���v�į��i� �_��F�c��;c/�CM�9bף�uE�%A �kpif�1��@X>�����M��C�c!1C<I�)��ZL�oET�Y�"��YI�=+�Y��ɚ<�j�u@HC�����֎���L��)INxe�n�J�t�K58��Ǽx���13$�!��O���(&72^ůI�����|hJ[���!�`eY%��o���@��*��w%�� �Z���id��W�z���/$T2�k�6��A�J�ը�W jm�.P��B:��{J%��8zQC|���+�q`��~��,������#�,�2���c�7`��켇�F���֧4��I�!q�w�V��?��G<�Q�~B�`��j�'ﾵ��=���@a+0g�Aa�<�.,Km5@�pls�Su�5�ra�ôW»;T����U^��o�:����c�%���g~��|}n��G�G���N4,L\]��}9����6A�� �B`��臽�|��{���g����Ï��Z���Ѿ�h9�j6�y�`C20#r<v��;<p�'6X7� :5��8+
D�l�"�9���>�"o���5���9���i0�
����߳h�! ����"+N��"me��:Ք��a視�%.�����7C~n+���/�Q�$�j�3I?�c��Z2g�ck�8��̂��6|W���	���C�ɡz���)�Aq���H\��#$MN���v<0�u��rOam��>�����\L0pb>q��´9�حݥ�9ZH�]���s3'�_�"ʯs��\���.��7��n�B��������o��6����M0J� �W�A�f~ԡ��6
;�ǎ�C��u�'eۧ7I�]��Sx�K_h�;O���VΧi�W�M3�L���?(3�9�ľN��.�LJ��E�R��9]	e\gg6��^���_�����n�0��w����[%������7dn��ۑ����.Uw��NE;�_IK��0(&��'Q۶�2�h��c4�d\��:���g!k \�K{�D}l� �Bߊ��)P����E*�֒������bˇ��1܇�/������h��4���PIr�:ڃ�?1�vj��'�F��p륿���p�ٴ��1�SQ��K����N�i}rr�wǅ}�'�C7���/H�%.ޖ �.�_����ݢ���V���Sf@����?��6V�E�?2V������꩷���P^�u�S.�C�^�3��,�r8H8Qדs�V���m# �����5L���(+Hl�l5y���s֮�'1=A�%T�F6�x��4:hw`�JzaU�����g��Mں�^c�v�^�
s���d����q�b��4��c��3ő?6vF�|H�7�sw���B}6�ۿv�P�NA�?꿁mB�u��cڂ&7�dL����ί��u�A�c MW�>�;B���9���P�b�AH?p���c�8G�ns�C�>r�Ҍ�p���M&�+��9�'���KBڃ5�J�BE��X�&])�E�Ɨ.�0��S��V�@|ӵ�bhj�sF,�$��z!D���@IB�*��k��Xӏ���4OW��CL"��������]6N U���+���Kx�يD��~cN�ui1�y�l����8UI|�]܊P��aϮZ���R�Fg���\K]e/'���m�O*Ga"<}Q=�(�m���6~�|n+����1e_lF���4O�s.V�R�m]���N����z;<����̧1�ۙ�%$3���Ntd�(�-�!�V���=P[��a�2^O�1�,��/#�κ�u�A��?C����=-��?<�x_���z�eTF����	����ĺ������!q�tV�`������Bp��������X��?��>]
b
���BP������G~�:w�.�_�<b/޴�N�	/��q����T)���c$ H�B|�_X�O�������^w��8w�]� C�Hd��+T ���1�������ȩ�|��U�x�rT�d�'�j�~����5U"���[���?���ɞtv*�oم(RZr���!2��p�N#|�s=�Ӳ�+>�_ �����"���ȫ�2B��9�R��j�8z
�`�=��e^.|�<2��U�&�Ԩ(宷�A��`V3K�l�V3ɥzض�?
A����Vf4��fї��k�Yy�>����wD�c��3�^/K#��^��=��F7�z?˺�m'쮚;=h���&=jy0b�� dN�\g�ǁ��A�ba
Hu�LNmt�o ��pD�����AҦ��Qr��rv��50^�i�(t6�s#U.�2��0�o�m|u6�=��j�Q�����Ӽ���G=4��d�
��4<
���,6��D��L$ق0)\���3�5{��)�R|����dx�[�S|+��0v��vW�A;���|���r��_��ۜ��w�$�͔۲�p�F<���U2
+�ͤ	.�[����I��?�[f"����x����m�؋/yqX#}����0KB�ϫ���Fu�`<:_5D5
��y����=f��M�~��ѭ���툻��U\�љ{��50c�w�����[�o����d��vLh[��Ƒ%��ץq��l��`J=&�)4�!	v�>̿��լ�ւ�x�������2��}I�}LV<M��S���W�>	� ��>�k��?�z�3��g��E��d��啲5"!�N�`��!�v�/�9̤4t�;"J��u�/�1ٽL�$�>�k�b�#��GO0�M?�-I����t�!�I���gu
b�r�7�M��Ll��,`�z'�Q �hP��J!A8�y�i횷@@�5e�?�-�X�G�G��C}���흲"4�5��H�&�