XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��s����
.5���'���S�2���Pe��rLN� >�) �@�R��>Uv*5kNP�����m��'��_�����IzG��r���\��h�vI��i�s�J0��%��G�P�u�~H�À=��w�\��}������:�� ���!��9���t�/�oീ�sӓ�Au7 M��V�P�4;y#���ȋ{d���;��Y�����Ck3�O迤-ˬ�}b=w���^0���Qa���uxi+�۰��9Њ&���B�&ѤY�S�5OZ�z�+f+�;�N�:�$~�V�B�[Y��ݮh�tϮ<1�a�ӇG��m'�a]p��.�Bb"Y�?�a��'���z^��Y�)�==��z�:4�1K�
��}S�:7#� Z��<��3_���[N^�s��� ���&�CI�}�0�^�PE�u�`<�kS5Jz��Y�c�\�lj�C|/}�~i9�!��%��%`��n��N�?�l�G/���Q/.�%�5�vH�Ϣ��R$��LCo�ݿ�HZ������]�w~T�����<�RbD3��>�^����!7r���cǸ6��zܕ ��F��~�{@?����W�k�T��ff�LG�(�~��m�B �\,�����&+��2����j�$����I��V��G�������� ���¶���[�%|'�0J��*p+�{KC�>N+lX�X�`�vr�	�R�����K���.& ������k�����&��	 XlxVHYEB    4013    1050�lVxI�ğ�~�gQ�i��ŲX�w�a�`�pL�u�J<b������lb�H��4z�^�ʌ�T�A�-�~��񜮡�����-�C�O�I�@m�6#"�a����#�(;�eWQR6G�a5uNM(����xY�Ɍ����F*I�J�Xe �2�t�Z;=�&������������������u>����^���ƺ��Á���2%���7?Wd��-0����5�:4�H�(X��FE�u��
�݊C�spK
|2-���x���p���sG���7��������<�]ݲPۼ�����ˑw\#4:���P�f��N�'�����3�����+�󾍼G��P=b��X��y�8p��k~-�N7/�-K���44"5����2�Rh"u��
Cz���I�/���;��Km�;�;}]�V�X�ۙ��J[�P/{4|F#
�̦"��W7�W��tX����NJ?a_�&
07��G'C�Nh���<�ro<���4���9[�݅\�-�^[D��s�qa��Z��`��=mϸۼ}�6��� �
�Q#/�y����;�<�jH��W��7�yo�{���Mo�>�t���!�b���FX�~�lߥ��}���e�T�}q��%a,�6-V���TL�]] 
;�uLܛ�RV����k����G�W�j�(:���H��ҩB��X�f
ӪD=�Y58�"''/��: ƿF!a �Z-�������x4%��.��8�������Z���뭤�/@(����#gR��u�Uʉ��J�,�r�.�R�% %�Y�Q�La�EG�sQ�/[��6U�bC�줷5x���\$���D�*߼<��ذ����D�J�Dq�A7xΙ		������fa��s��߉����>\D��Ĩ�$�r������
n�]�?W
A�ϊ
�ޙ�=��j(���2I�[L�.b��`��jt:�]V�"ϒ��L#p���Zm5�:i|0��.�De!s����c:C�/f�u�yjGաi�ݤ|��	�G_�G
����X��E8�b�K�#+|t�=�c@	�x��,	|���p�|v��a07���)�g� �~*�X{�"c%�#BkiG  ��r#v(j ���N��������Ч_�sM��]r݅����`
Rכ�ձ�T\�Eץ9�6�)�ҝ�/0z?��B�ʫԃ]`�
˶�%	�(7�u��G��j��8�,;3�4�理�[?�R� �����m_���T��W��\��b��P�E�x��� ���C��a�`�;_����B���q=�`>��"R�b1�7&�R�a �Zzq�$n�ˑ��v�J��14w�%@�}k�H�Fذ�;m�:b�U���Qk�=�p�t7_�de��v�\8�N�]�@����������l�4<f�B�� �P(��+�:u�
�;]��L�b+;�w���oߛLP�s5���U�6��5g\�?QPD��2_-��>��e����f)���֒����u����q���顲G�|"�&���]GL4q��:�m�[b2��Z��>{S��%:ϫܐ�� 0��F�S���!=cD�Q�`�Z�^��t�����C�Z��).��nB��?c�c�Õ,9u�P��ˌZ���� ��o'��W�'^/�������VN�A�u�2J.%�&X������Q��{;A����
Q�mĦҮ�]mT*R^�]{ύ�)��W\9�>F[t�;����w�<(0��Qg��oޭ��_|�j�~n�TW멲��N����{e�ҠQ0ET�P�a�u��8��h�=�$�p �`+��'jh�nq��*O>��,����E�+���)������)؜[�"�%��Q��j�ĸ0�8��>|il���;Gb�i�㎉hi~EVm���?��N��|%��G�9`��t�n�T3�ѿ�I� zcRx䚽�㯜�e�d!�a琍ɥ�c���ERcL��`$�ųYO��
"E�I	/��A���p A��Gr[���mmqΜ'��)���Վy�I�g<�|լ��Mb5�<�<���W��y�r:{���<f������|�:.#����_��~6��d�y~��(��Щ` �[�	Տi��>�:�l�
j�U�$+�����a�s���V�����X�M�I�D4~�]�� �w�F$>D-�`	�E���lp��$W�uh�]�͕Fַ�c{5��z2�T�_s�%٥_ �����l��:�$(���)��G�V�� ��2���?�Ƭ�$�<ѥ���MS�A"T��X�LT��8F�Փ�Z��/i9��)A�0��Oc �f���j�KزT���a:�M�%A/_��j�!�"��F�{5(p�i���G@��9HR�h��;���,{|ĳ��A6�ʲ1z;XrW � �k�A`j���[�NpY-s�
.(���~�ɼ�q}(��%�p�o"_�N�����-�d#)\��9�����#�٨�N�]Œ���/|�����b�k�z��2�>�t��i���-"�������M8˥�mB�2̋6��x�x脵Ew���+���(j�o�6���,�njbг���:�
�uՊ�?����J�E�=8��u/�G.�?b�w����U�A9z�V,M��]P��{B�$F5������#>���"��A" �A+�~PvIbR�*�8J4�9��#����.Dx�lr���*n�h�����,?߯�e��R�=f)S\���d�d �ڸ��b|�����%��.��l�s��pӒ�]�����kO��-(���'_Tϡ{��
;)(������M��פVgǧ���0���'�S�=�^��8}���R��s5Qq��>�j����}7�1x���ɀ�H�l�G� x�Vy=h�L��[5g�?�}=?�)�C���ìjD(WaU�;�׆���r����*�P��#Q�8b���eb��4���u�<ٕ�<�� q�}q�!�ϩ-��9f�Xɳ�ӏ���
�r6{y�A�����<͝PL(�Q	�~����cu	��f���� � �YW�,	��F;ì^8j�������b\%��� ���� 1�8��>�4~�[�L)HNc�_X�z���w�H?s��+�S�;�H�l��u�T!�-����3NkZ��՝�e$U�աw1�8��k� Fm�y ��VL�����Ӆ�B.�-�LȺ¾�"H	�w�)����W)��]P-X�7M*�Ĉ�ii��Im����x�������m0�U��P�{�S�`����W=0�(�U˗t�\+�ޡjh�{�_$f������񊅶�٦�Q�]�����>-Y�5ǯu}|~$R6
_�\ؒ����^�\2��8��P���#p�Gg�)��S$El)�JF�2w���K&� ��l�7���Z&1�c��
p��b' F��E��y�U�"�'�(f �5�����u&���)�W
C@>���]a���ȡ���xih4e����f��{�}C�O�?k��{5g�ߎ)4�7�uG<SfYiv^��B�-Ս�b$��ٳі�� 4��R��ͼDLM�#	L/��%eB<��
:[�H��׻�>TG��wi��q��Le��Y�fβ�^V�8i'�\Q����_���[_��B�LԬR�4���c]�(p��-`��
ۺ�e�T�Q>��^�5(l5�c9^@
n2�ܨ��xb�^��b<�1
��_Wոe��&�AI޵���$�k�����Y�o.qw�
N��q�I:��S��WM���潁RuK3�q�T n�ʫ�Z�6R��(��������G\�l��zr�]S7c�#�Gr{PM�����-�2������j�j�:���n���t�À�)/��4����^<�*O�^g*��5Bo=/i>n�B@���	Z�|�S���op��=i��Y|i�Q��n|���3$G����3#t���a6֣<F��CN0C6�Ø�3��@<��H-w���D����s�5�8ګE��+�D��O(�M͎3�+��f'��Y+�첹3��v�F+���.؊���}��F5n��R<��/�S��(���/8>eu�{�Ѥ�+���\k��P�
��sEٝ&�[>Q��"+RZ�YE;���O�