XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��
��+U�ण$��"n�����m�?���?��R���&\�H���]�Ê�������9d�n��n-��\ڷ>z����W�M�O���e ��?��ɒ��d2�p�
W>䲂���	N�en(z��͌grt<��
�*�{��~b�6m؛��z�Z Q8���%YF=�y5`��x�ĢS�0���p�0>�e>�M�[�q҉�����V&L��������0ɝ<���vN���7�lu��R�����N��-e6���	,5��'m,��/bs��禆�����W��eu6�Cɠ���ю/��5��k�� \��&'�R�)�֧��r� ��Z��C�����E�k���a�~|���������mS�����Lc�����1��V	���'}ā��Y$�P?Μ���
演���������dKX&U�0Y�|�����![e2_\_A�����cn������:5���J6&A��]fI�g���m�q�]�㏉ɲp4��ÛmE՜qk¤�A�j��GE;���q������~~�A�J�l4X�1���Y:�XW�%]W�ua [���A�ɧ�����XGA�b�c���zN���;/])%"�2����� �h�&�<Tf@�J�s��7�|�c��T��7�)��4*
T��S��o��?�
�����A�9u�b����-ehY�@�K3v�a����'�j>����p=5;R����$�A�1O��]&�{�n~̆�$�#����H|�XlxVHYEB    3189     890C�?V���.}�Y�Ag��v���4�:��T4N���zk��1q�a!@d��Z�����h�kV�/t������}eck��E����7}ȩ`��C��}W ��a�Ly����!��vo��k¯�l�ӛIM��v*!��Wx4�y���yS*��M�ʫ��  A����|��T-X�'t�B�%D�o�=��w�ߣ��|��舐e��Ɣ�ϐ�x����uD��Δ,1א:�Z�_\|G3��"�F?��8}���5sdϚ^k��y���ق�m�,Ao�b��H���y�F���vf�L�2�v����X�̳[����5O�j�(�K"���gz�{�f�G2�1��*T����gײ4������0��y#C���:���nH�r��+IT�5b��S�k��*�,s�^�4��������j�#���3��Θ�6MZ�%6b,H�lu�v��RJ�<�$�V���`K�b�\���麵�_�w"����P��ں΃d�E�e^��0N�G�,M��mD����R:V���.�Ij��iٲ�kƭ~yת�o��	
5�X�r��# �Á/�n#O���U�����}Vm�3ʱtc���F�S�2s�<�H�a�1z�n��2C/M�vM��2j�Y,8�ox��':��-�icsQ��2ۅu��2n��M����{�g�� g�m;kе��\t��ƞ���.�p���K��k�Q�XՇ����n|b�W{���x7���\�Ѿh�ULy����P��g|��BgI��i�$��߄�,�W<�D�^raCT��e:8I���^߂��դRJ/����H��R�T����t���Lu.lwjN|�-�v���z���͆Ā1�^t*�Y)s!]�6�@�XH�f���g�y3��L�2,���bS*�*�� %O>�[D�z��r	��W����2�E��ЃZ�l(/P<d�a��E��VY�u�����������8`���r"��-JM
�'�l| ��ڸyǙW���u���3���(�EK�2��Gn��UqN+\:�2�@ �^�n��AN�(�3j����_�C�d�\�X�����1�o^.h�Fb���'����D���.�G���Һ�z���4���[1��YH�QY�p�)n^B���1{����gn�Q|�<�O���u��́�G�A7Xq���p��5ޏ W�:�'��!�>�Kb`��Er� �>!ujs.��]=���|�F������N=<	6�u�6c��nn��5�[�ƅ$y���x6�@��Vԧ|�k���?�((~��+�u
d.�O6�U�9X6l�i�7��ƈ�Cb��[Y�B���HlȬJ_F�U�n����e�4��oP��:6�>P\�gg��j_L~x�hm�\s���	�'^��<�{��J��g��?9^�t�iջGe!��ۃZZg�֖%:���*g,�}��W����Wv�%��Z�9�t����f�j��S��G�������X>��H#���`�5J��"�i5��Ms�WC�n��m��t0����|����Q�(���ԇ�~5�����^��C����o�χwR�&'i�Ʀ?��.?xi_=�C	���X�'y��䡭1����%�k��#�x�(Y�c��P���\Yo��u����v|m��Z��q(�OԣA���M���v:m�������R,��HeXL'���k�ISnX����a�%�҃{g����r������^�PvES��&��c�E����c�·Z��85DUc�>�����G�H��
�_��9lƯ����`]��W��<�gD�L����Pv6:��}dmZ�>k���l@�;3��R�lAܴ�#��O�qF�vk�ALXmH�(u�'��O��Z50�n���1�ѥK�"d�
6DSG�HF�b�3�M������CrA�W��N�}��	i
HX W$����_#�Z�_0�-��̱��WL��c�;eK�ř��[�]��O6�:3Ƕ��|*n��N�p���K��Ş��#���V�KZk M�⨪Q�7yY=�l6-u�x��4&��_5a�?$��hC��v����e��\��M8�!��QT�&�� �P�Iqn�2[3!z-Q��o����C]�J���R'�bk�h�{����[%