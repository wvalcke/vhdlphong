XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��T���= eoN�b��X.�;�X�!�PW��*p5�T|�1�+���c���70%�ha��B���@������DIW�t	,#��K��Q������| ��ԅ]��$d �#_/����i@��K��	S�۵sʮ�Ա���p��Gpy�SL #1>g.ג�4V�'�}��Mb � �Q�K;��.J��� �LW��K[a��(�Nf!�����Z;�<��$E�<��X��-�����d2^��s�`"3y�G������%Fv����C^�ִlZA�5Ј�<��AVnw���[��9?h���	�=V�V���	m�<���O�*L�7�û�A���UE�KtP�6�#�����'��Х���!&�b�܀X��,đ�A�:+���G�ʅ�p�y�+��:���ti��Hz��Ŝfq�!fr�'A��h?*Ƒ%�� ��v�*�!�jU�{�W���3��B�Z�{���u����bwvA�ׅ�p��U����Y줨�BSs+�ܓ%]���or�uEY� �<}� ��K^���5��	��h��t��$�M
�!��ʝ��R�sNg6�J��tL'������A;�_�"��nwr��ʁ��h�Gw���}���!�`��Ar��b����H��Ν� _��ZtШ��Z��!e~Y�����4u��۟��Ť���y7�z�N(�U�ɀ�(&�/���C����qܐ���C,��u�R˴ �Q*�'+�XlxVHYEB    3357     c80g�[X:��~��\	>��dg�`�]F�\�?�A&��o�����z��Q��|l�_�/�NN���
�n���
 ,Ϗ��6o�$��*�Q莠��5৖�D ��D�.��L�eQ"��ã�aF��{�f���r�1��r�½�����G1$\<�� P/!TS]l��!�bU��y�<b�1bF��bA�,l�x��)?<9"�۵�a�w%�ϫ<����;ǭ�u�]���泩'�j�U&����K��H��sd�M�d�b�X��	�{Tk)����b*���My���_3c#�ʇ	�U<�B��LZ��&K�8��@ т&�lf�f��j���K����@�x8@�w��/�xLӂ�f�ͬ�w�=�(È����-��"���7`I#�y�J&�4Þ����TH=Cn�J���6�] D��U+ZD�.��� ��BxsRi�< =�5_j�'�$�B�%V�X��}W7�����8�A�	;�~�DC�lFeU�Ҥy/[Wa"�8�bs6Mv�)�,��ǔj��Yep��.'T�P<a����p�=l7�1��R�)�A����o�G��+H|�M��#3���(��@l�s��Hc%�D '�r��Ƌ���9�ug��
�=՗h���@݄~��IڼIU\P�r�c$u"�,�w����׉�}�%4@���!�gj���u�TF,0ȥCޕ������8&QQ,-[j�H�q=;�l�=��7�d�� �:�}��\JehZhlzc{��0���Gx��o�}!����x�q�h��L;ʽ���d�%���*�G�����ޜ�Z��o�d4�ra�n��8-	��ռB�j���:���-e��rϛB16���1:{;z6��!6K�e������s�Қc�O�V�SKRL1A�{N��zG*��hK�J�SHfOr�K�l��6�l*�Lo]TJ��I+q*��Q�^�'��T�pY�S�q �|�HY�G�'^[����:)P��V@э�*�h�{�7�3+�
h2<��s��"�v&�b��=vX��^�l-X���1EaͰ�TzF�;7W�t�am����4�X_��*�z��.�*�{�#�А���l����w hq�z����DVc�y �4z��Fg�.�?;<Ќu�X3~�$�o>�qeMԚ
p��4�E}; .T�X\���`�YA�m�����c���iz)[N�uq�"�n9��mv\G��/R�v�UP>_��m��~=�����fBc,2��@lvyժ q4���a��&c�6-�����C�\����R�� ��C�T���x���s�}�ց�u�����USN"x�B,qGE�W>��y ѝ�sM���T����d_C��޶�;I����v��b=�Q��#�V���]IU�^:ym�82hj�t�#g:������VNE���s�!�ߝ<��|�NO��lRA���#q�A�'���S����R��d�qM0����[� �y<�6����t���&v������b�e�5�(�P��kF��|�MJ�iX��6��ّ��]�)Cؗ�y�G����R,V<�H�>�Pڦbn�ɗ��k���}�f�D����y`�?��Z��z���d�5ȱ�Oxx;e���QTLjHh&5%0��~_?���'��:n��Ʀ\�V��/z�m��ٳ�J��M;&3㷞;4�`W����&\h�� �.;�6�ʗ�'�DL�x�H\��+�bk��q�R��x}�	�O�)^D#���v�o	��^	������^N����\b�ֳx�D��k�IzJK��Qd�����'/o�v��1wo&*6�71�~a�4� ٍ]���r�{
)�e�tQ��T�b�O��8�4�2�!���T��drd����v���q=����s���GzȱM�v����8�Y���rNIX�VƧf�ཱུ3��]�.�����>�H�Fh��R��.���V$Q��2��ap:ٷm�A�O��Oo�Zt�.N/(06	''��	�a��10W@��0E�t_k�Ê�q䁦�;q4��|~Z�;�m��!�[�h��g�]�)d���^&� ]�K:��3Yr`:�#Y�쩁��U�]iŢ�*6��)��I�_
1���(h�)T�g\��Q�{�|�I�:�4W_�$�j�M�v��T�gnΔpjS:*Z��]��������%>H�*�iy�r���a[�.M�ز�N��w�1���_����X?j�>ZR̮�������ț�=p1K�eE٦'=�x$0�$a?��6�NP�e�@P�M˶�������4K��C�}����VNV{Rq����eX�e2K��c��Bm�ym��ffg�B`��h�po��o�����/��G��9j��ee�HE\lp<�)@���8q1��qק]���4-�򭱁��Ů�g
�pK�����z��f�s	�>.��0��Y�S�a&�6�I�S�ϻ��|� �6��#h��w[H:_���W
�Fᗻ�KQ�zpb{'fX6 ��|0��|�"�`U�Hݡ,q>1P5���ٶ#g�	��α:0
��������$m�G��t��@R��v1��Ӟ�0��d�r� �#��,��lz�z@�N�Z�s(�B�s7&�n1uirR��"!֧��4�=�������Ũ��Ͽ߇]�kla"�(�cY*�K�
��5����;b�>6ɽX��̈%�|��]{�A։j�S�iG:�9��0��bT|O��*���O�Z9�����B�&T����n_��������4������(̦OWF�Z1�%`�:'b��]ۺQJH�VbX�U�јa���2Z�h��I-`�ʔ��O����B��U��%Y�
)��Z��+o7�)�ϸ�UN�(�|jDZ+z����i��=����NI�r�"��+E�<����Uf��W�BN{�!6H�:1�<�#f�X�vC���1$q���X�sgw�By������9�lƞ��R>�n���7����/��1�(�2�I�
�V��rV��q7PO@�:�Z&�n��Kܸ!��J��G�[��7��#���9HDd(��߅1O�k�KZ63� �,tw @a����b~��*o�%e]�MZU�E1\��.���N�z�F�H����ݯ_H�f*`MK�&����P��