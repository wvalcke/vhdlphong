XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��P�F؝�����R�?����H�%��s!��$f*��>6gl8[�vqh/���z��Qw�,�r��Gq.��~Ts�C��],g��ۮL$�Mr},�@Q�C�*�8�B�:�!��{�%W�d���D~���*�%�qD�@���opz�s����\����k�'z;�Ş�]W�O�w;�wr<�E�Z��"�R���-)<REw��k_�0����H)�����m/���D��"�/֔��jp�`c�(ƛ�� fN�e��_t�w�w4k%&� �K�P6�����Hl��6$�[f���;��߼�W(M���+�,�V�<ٛ��n���lٷ��*�n����j���;����=O��ǥg�0���"��^E�m���'����>�?�@�>�ʻ�M49f��.6n�s���q�6��Kf*�w��]�;eK�{�QH�)��G�ԉ��"+�E��r>�;����x��A���b\(Q����^+T�Y��O��2��K<�Vh��t��!.&���o�wf9^u�JˬR�	��X9H3q\�Z��P�b:�HZ��9�M�oo}��'��WP��r�������	�M�å�+a_���$��ww���v~��J�B��	�#u�'j;7�:��i���H�����Ȟ���	���^ךٽE��&JO��ч�t2�&鳫�ZR��B���a��|F`� �]rF��F��{!2S~�_����Z�`ax��>5�㽚�';�bT��y�%Q&�<8�w/MXlxVHYEB    6e28    1620� L���U���XwS�}�Ɛ6���� ���|����#��!��$,�eN�^��A�I	�.��ľ�]0/I���FK�����(�Q��q�_L�H�92Hu�$�Y<�Op�08�rW��I=�V�31��=����*��°Jl-~%<e�?��T��Bk:Yct�^�>Ѭ�.\�y�#��T/[��MJ��`�]��6E��9>ܝ�Ͼ��F眒�s��/�-���60��2 �dC0�/��O3�^�h#�cB�W�~+�3��Hp�e1{�"�����s�<+@�Ѫm*�({`���m*{����W�=�f�5���	�s�������@��j���,540,�4�/_�)+�\���}.()�p��������jv8���/���;-�=}�K��9)��W|{�i��k+�\Td8MZp�5�ez�C���kp�MՖh���ў�/&����D_��=�4�]��}��{��5�����F☣�tN�Qt ���������J:�P��_3[�F�G��G�-Ys�d�7�{S�d ��*�Y,k����U��w ��M���ՙ���Wݿ���#	�J�?���?*SH���|֛��G^��,�麿�7���ԡW��*օpN�"6�?�ʎb�`�tTF#��3�x��?w���0
��ݑJ�h��mV>׾O�Έ�����h暎�f�u���<�bR�ߦU�ӱ�>C
Y�?]%�;Ե�,k��۾r�aR�� +�w�ü�Q�U�]\U�J3g�DF>�����WG^/d+��Uj�ѽ���y �!(�P#������p����k�Ш(��;R�E�K[$�k���z#E��D�Ƿ��%+���m�x����ˠ�=�i�^Q���̩6�I����3B&���y9���"�٘ ���T<���LV9)�y���Xy��Vt��~-���E��)1D�{d�'N�.�Ǧ��z?Է�/�J��W��Ʋ�W�b����Na��8�I��f������{Z�H��\S�<U�hM��ʃ��w��Dy�2*jt2�=t���f���d'~#�L�(��^Q#_$�ב?������%�f�hT� k���S-��w�I}P(��!_F��ԩ�q4b���)���1����M2s����I-I�NU�!��hG���#B��8�����_���� �o�M��Z|،�M	د��t�ǰ���R2�ä���gP8#�{/4��q�kq,�ߛ��{o� �c[���i�И7�)JZ7��?��X���hb�u�]숔V^Z1�(��ȗ���W���țռ҈T��=qv(�r�,�笄����~kYTB���Z����I]*-;v���r��o�|�ȗ�Rt�rm����{�)���
z5�	��;g�q����ӓJ�B����Di	��R�Y��쬁����\�c �+����H�0 O�|#k �h
"�2e�/&t���8u\�(��bU���@�@_����|3�,|�]:<}A��@;������>��SWo9#���f����3a��2���JN`�jS�sP���h�����Ί�/O�U��g���;چ�4��wO&F�j'm��)Kl��b�-:�z���M��O��>��=<{���@��+sl�!�S�3RL��P�Av~��a��k�̲���� )�բ�b���.;Ğzz��(�W�㺳���8PJ8܆���|
�9t�����GϦhˁF4�NTD`m��/�{Ae<�e�{�p��(�t��*~u�e��S���o��L?���썌O���,��K��KˬQ:j���)�G~�s��1�b7i9��I����Z�Sa���
�ٹ�[��d��N=�3�u@G0�:!H�Re~�x��:���D�9�"�_L���7��U����� ���3�-
�Hc���<��\D�145�	X�F} �^|ݪ*F�*��I~2�P+�� ������r�l޼��@�0=�v���'e�����n�������C0��09�3�A�;_����|¶Lo�ʗi�����������s�a�tb��}` B*��b�xR�zL(�`.��ܥ��e�O//���W�21�L�����	[ͅgce�����:
���a�G�Y�e�I&���F������lkeǁ��?��܌������p#^�A3�vDe
ձG�eNaY5��g���Y�uu�������j�(����'pد1er�QL}R�.r1_t=6� ��A�{�#��!��������X'��/U5I���Y:�xfDnP�w^��J)����Ӝ Α��e��%|�~!#��O�ԱF.8��d�F'J�K�x��q����4������K"�fV����e���������j,&��-[I!
��q}IRBp3���j�o9	���
��-���1�:~�ʱ�P�ҫL�О�Uv��Y�ݳ]�2y�g{�!�g�oo7E"]���qu����Ƨg��uP��x�
��
5�m�OU��R��Ҵ�eȳ�(�S����3,��B�0�\���X��%L3(�&�7w�Ӹ�C��D�}Ɠn�?$�h~R�Ҍ��lP�H��.@�H}��ſ���){�V�C�$c���%q}�l�k�o�&nn�h�欏����	��g�N]J��hH0pk�!�H�-O��F�.U�AB�x%ȍt�;���JL���C�7����7`��/~75+ �<q>m���t_7��}Ey��Ԋ���mr�Uz��<�L�8��Z�K78� ��]O)Y�	�� ʃE�c��A(X��ˊ�X0nD@������G��_�6�e�Z���xw��b�:��PJ�H�ҷQ��r�Ѵ���l}P�㻑
����>���Hb��AA �	*ɓ����kėr7�y�p��"�En��C����ɣ�K���?��u!x�Ƃt]7>�2�i�k��5~�@�uo��O5',�ڪUlIYa
o�f>���4���.��+�Q�a��"�4�چ�B�[����!szΰ.����xD�����ו]�A�8��]�g�bQ\\�x�xF:p!~i�o{��:⭆�Z|�]��M�()��Lg�E;p�� �������BH���-}�`�)g4B(�-Q=[��՚)���Wo9��
nߺ�����KXk�AV����9���`�O�a��]���M��ɲ�c���t; c���*;O̫��A	�A�a�ɳH��ޜ�l���(כ�����l��\�F������iq��h�m\�MvZ�/|��=�hَ"���C�(��0wδ=@$�+�jP�Ne_ծ���6�BM���TB(���m���XN��4ݒ �g�]Bi���^���8`ZY	��?*bu��vDں�IP`�n��\���
q�e�sL���r� 0�Jt3W������8���l��J���7��J��`h���BDMZDX��əq�
�GL2�p�$����lE1�&�Ԙ1S�� �wtA�#�X������LeΗ���%GӝK\�1����Q�j�qlqİ�$�+�Sc�m�+�MR�ji<�*��;(n�X�Y�M�|R���kg��{eA����L/�6����4��đ�x }�$�$�aL��u�S�/P��kԘ��]�<�����`��8���v��5��! <�%���&|-�yuI�����;#���*˅f��,T�Z�]ٶE㥣�Ww8~�{�6���?ϒo����0�Z�in>��gR�/���cn$����$�~^������&S�^h'�j�\�3�[����CM3�ʽS�Y���Y���J��|�HM�W�yf����h
Pڠ�_���|�������>������&�B������	<t���a.�[9K*bW>�j#�Ro9�;KP�3��"-�
6���G,o~,t?i�	����tE�� I�^Ű��T��M���Q�䢕�ʸ�};���u����-0��9�U��_��h��}����(_�Z��G(�/����.�bn�ɘ�0��ߧ���v�e`|$j���}T���b��c�%�|-��M��j��K(�$2N�"�戌Y�H�џ`����~������=���O�!�E/I�zPO��$�FA�p�Ҋ��8P�rr2?��'I�lSȦ�����ߧ�BI��}$ޛ�������ȡ�35%��[�� 7$۵#�y�$�@d2��`/�f7$O�@5�2[%PQ�s�^�y:�p�	���M�@����@�)��؜*���:|��{qź�9�v���^�ed��̺�n��+�����?|Q�ݸ��&���DU�	��ʑq]� .�)Y��Y*��}S(�$&4�9��X�D�G���ұ�R����x��IB�LV�M�#ί��g
�dTܞI��`ŀ���<hs�J���ʘD���
�jW�py�LPVa�+�P�s��������+�0"�T��������=��A�y�E�v�,������*�XiAa���/���>��܉��Y5Ǥ��D;�� �-�aZ�ːX��μ�'[��t�	ԌLr�bmgw��t:-���8�<6���y�{�Z�͘��X�Y�l;���/d�z��_���XF�D�z�%��g�ScA{��?m��t�z(��.�[���8���Ot9+6F^E+L��T������k�Ok:���������g�&��݊���X]}܆Q/]�-؆����������e�φ��V�^�4}�ĵ�E%{�BhB�9�=�Z�P1�ȖuB�C��<��F:�wg��I#�Y�v��g�4}r^6,��񘂿n ����q�ڋϚAb�6_������1"���3��Ј߸��<���xp�(�Y�@p7�8����Bʇ'S'�����xзc�O����NV��3��A��wj|NY2ЂWA�Z�j�6W�ߓ�5�3{+BGZ�I��x&K�����#���3 ��y�/�\�o+�!�{>���+C�~�#���ȫa`:�m+"��)ɱH̓���o�&[��]�Pq�Z)K����覥�ޮ����(#5'�[4����b8��Ib�%�4�����V �Wd�I���bt�o��Ngc��6&�^3;Xl�_Ǽ������L@����P,vT�܆�;e�N5iZ�x	j�UQ������5�z6E�J���d&R�R&���K)s�;��y[����oW7c��G��0�����9r�5	C$��9'@X��MM���B	��Ti������6�cC����4Xm	��Z��ة|�ǤH �C���ի!V�&��/?q�~��aS�#:x�k
��P����ں�5cQ��������]Zh��r��E^#�"���U/��+��0Y�d������P>��3d�y�)ZP��"�޻WD�'�����Q�3����?~&��s0����#���1Fl�m��Sӟ�?��Y���{b���֓վ�X﷔��ed�ĳ��T�F�C���Q)!|�F��>��hk%)����;�D[��X��j�A?�N�8�%����)�y��1�T���