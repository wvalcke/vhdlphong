XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� �pR�5Շ��2 K2@��;��ܽ���T��6���,�*��;�֝�ӿ]��ć|)�S�����%�� �C����1��4Q]�o���s�h�>ǥ3位@-�Z�tzPr?e�"����6x�^K�G�c�X���� �U#q�b��5͎������Z)�����V��Z�����Dg�	+�@���L=|�lGf�}�'U�Sb<t�瀵@�:��q=���R`p๮�A�T�0���eXTsm����K�?�=�����y^RBBB�cI|�+�w� �=03FΠ���V�Yl����0��&>^�Z��+���;w���ŧ�A���&;�Ut�'��ь�0�P�i�s���OW���NM�����y��K<_�ՇL^8|� �`�VF6`Xf�{fiE@��G���=�o_?�4T�e7����c���6�F�q�@�7Q*�v�k�{Qh��Un����M T��g��\������7���z[��2��}Ǽ��8��&�+�*.��C)�����P�{��4�+2�X|��n��V�Vߚ;��t��<�!�auɴ��%�G��E�2gc��d�w� �hR����4?[�����9�ԉ��a�-"K�����qRD,=b%��2{(�o��e�'(w�&2G���B0ܒ ���n���D��� n�$yJ���kѱ�W�Q@����Ҳ��d�-�1�q�u;U�d�@� ۑ&��̖"}p���{4��-QY�jJ�T��]_f\w��	���A̮Ɛ��wBc��XlxVHYEB    3d5b    11c0�g ��K�-�^s#;�+VF�����<eU�n}�?&= ϼ�;$[͹�Ӆ���(��D<^ǚ��s��yݣ́`��R���PW1��S�t^��~=�"�vW����0�#�V
��:�R�]d!�>�M�����[���u5�4:5��F�`9��5���]&��w7��� �<"#BxY$��L�_y�>=w�з����YVG�G#qz��sYT����.�{,o�W�P�k�|Q����e��+Ӗ�2�ZQ �����p�e0�V�/�v�28��疷�7R	�%|AѨ�c����Mo��Bױy*�I��B�����j��P����1l8��v7�z_�\�3��=��x-��ny�L�$�ni�3�b�=��,�O���޽�\���Þ�w�qT�Vq���b��!F\8�*X����Q9򆃀�$��i��k����؝b�(%�Kg��Q�)�Gj�u��h�4�F�K��6�!��ݦd�H����d.��mz���-����$_��7��eh�� :"R�������`��f	:�����Z9�p^ymLu7�e���㋼�m>P!��N���*��28�2�*�'Jb�����F��IE 4T��X�Z
�r�Rf���@n��M�*�ճD���%��h9}iD閖K�k����z��k��=A''rylbʛn��9���s6:��u��LU9
R%��}H`����t�tf�>$�X3^��uퟁR�.v�Wi4��w��s�j	����<��T��@�$�v�)~7I7�/��L�^~��H�$
	]?�aX�i�\�m݇F�UrK��
�%-��69��k����+]��~�\����
�tDQ(���g��@෨e�}�J���He�T�]�N����I~
⊩Y Z�C!m�p	e��{VQ2��a3�W�MQ�L��pԕ�?W���9�~���h�X�����IpɽP=~�Ac�B�q�\�||��R�.�sݺ�������
��8����:����|�c�,-̳#���B_��/
�_v��#F��Y���s[mXfّ�S=��f'm����p2�Pp��?�P�ow����b�������o�&C��tA<�ң���h�1���Wh��Cf��f����Fr4?��ye�:&YF�����G�[Q���y�ZK]��W�
Q���Ѫ�3��|+4G=F�+����[f��f��o}����G_Π�=�4�1�d�ZBi�s@�P^X�$4U�&���=��8}��!S�|��ؽ�2��㸏F���x�Z������H~[l�2/��}eͰH4��~k3�1x��_ɇgt%��h�"�bAs�z�=&!eC�А���ws�>Y��鱁�zi����'tn�,訁��h���F��Drb!�@4��H�cp��)���{�����l�zhxơ%$D�_��D,�׼�K�M�B2z#�׭��Tv�����2|J�^����h`�^���*Y*��a����S�FK 3q�����m�hTt�Z� �C��[I#���\�_��)�Fv�
��^R�-���m~���83��{[����=�W����D��C�m�w����>��zQj��D=,^�٩�>�C����,`�R���ɨK^�����7�r�^	̾k1��!UB7�x~K�� +�ښ�A��u�����ઔ8⡸�G�%�V��?a��߇�B��6k�>Õ�"��wj3)F�E�2�M�?�|ҨM���@].n���)�u9���{���fIݻ��������4_ �t����9J��˅']�ā���5�v��%��G���eޖ�i��z>;���H�n+�x��,�SY�/������wӒZ��H��e~>D;��~��ș�Ҩ9g��7��ۥD���%���tq*�pyos[�@�g�Q(�~�G&��H��+&�}������۾i*�3�0C��c���昈?ؼ,���6 �������[�D�.�=�ςS��ӱ��4¡����"�"���H�DQQ�j���X��jcJOO+�Y�3���ṭ�=m�J���d��;D��z�>$k�l(�����������/}����W�6m��5-!=��֖��1���G�#�����G�y�VD�.�X+Ͻ{TB�KM��?:�QA�?[Rٿ�S�i���Ҵ���<'`�[8([��i��I �lW��3�gk)I���/�+�eU{44�/^(�C�7���*�p��0Ik�:-�9j,������Iɱx�D�/��Z|�k�Y�'S�X̓���2��kC���X�C���<i���R�U��{gq���d>�1ߛs���#Z�_�6�>)���h�2ɠ�J���{F���r�[+Έ&��vܞ���a��,�W�q�\�$�Κ�ce�Q������@��pv"w	udB��Y��0��x �F1��9|�"hǼaeGҡH�~Y����:���H��xȈ5}��k�qwz剋��8�{� �a�X�q�:p�����\pZ�*w�Y�?�ve��`{E�[��Q��ˆ�T�e���8m6� ����Ͱ8ٌ�l�(�R��],��<���&WdA��>��]KB� eR���5'��D����8��ZNzu��sf���3w"!O4�^�,��zb�.G|�#n�|���eF��H$vWU�]cz����Ҡ�?~��s���۽�LHS�D2�d��;^��:ϑ�*�����O���Zk���K��"_��}�O��â�\����<�u3@����XXΒ�Ex!������ ���J���;����#X�����B�L�]�#xU(t_�՗z�T�)\�ڻ�L�5����ِgK6��Ӹ[��E&m���R3�����ד��D��<�.�֝ �Q��/��sT���L1lj28j��{�#4��f��#����C*5|�M�C�� PO[T��I�?����1 cE�q�跱�lU���A77���q�QI�G�0�l���m��a�2�Y�`��Y$n����d��|�7
8G����Y.��X������K�34:xw�;�@X#�e���i����C3?�Ѭ|
}��D>M����·�i���d�];'��Y�Y1��:�NsF��;Ps	��ƫ�co�MO�����;|l��������IRظ�R�:�ҍ��K�F��:y#�o�F�{�I ]�wk�*c@�=Α�D��KO���h!q0�t6־!���l,ae�(���^��z���;@���>e�����n���@<�(�>+�F��*���Y/˘}�R������Ɲ͒���m�b�����FH��	����bg4�v��	�`�>a�؄�B�Zw@U�]����7���vO[��2��!�hx��l~��w�p͗�U��p�@�%.�ԇ�k���W�[���Tf�o��/���IJ!u���ʓ=�Rʏ܈��0խ��� �ژFz��!�]ZB�}�l3`N�Ӕ�S��CZ
�M.�A�w������FҷL�ݬ�z) =G��������S�����/�`gJS�"�����f��*�1|��nIJ�O%�ؑ&�i��h�(3�o�C���O4��Z��ڍ�AfL^��~X��b_\ߧ	��n���P7}��"L>�d��+�~�*�(QQs�f���nqPc�0�,� ��u���0�u.�ޙQ����+\g��U��Q�2�_$UH��cUj���Z*e3�@rΡd{g�tXΦG�ڟg������M�'�� ��eq*�>�=ힹ�T:B�@fe(�G���z��!�9��x�cg �g�e�O1�m}9f)iCe޶�:O�F�B����  �w�r������޺��o�$���9#Z)������ٮ{3�<��Y2|k��r[���p߾���gL7�!TW�u��.]��^U���LC���жp��lGk��a�=��s/ �T�?m#��Xshv�j�k�&v�Y@�l�c��/F�;�v?ۚ"��u]D�=���v K����R*����w��;�z�h���z����9P(���6<4~&	=��B$o�*Z�P&�k�?q�<L|�S��B�?���� �懻Yl>eZ�%�L6��ρQ�S��p�����B�N�F�����qԳ��:M{F_��Q�5�I�6���1`���*����AV&���bk>4b�I���U�Pg2s�!uS�,�.���9Ԟ[Ծ� pY���@�j�o)��q�K�~�Ǟ�� }�%�&E��6�?2�ǞU�o&��-���/�=������\p�	����?�~@�L�N�^��xy��:Xɱ�!�$Λ�V������#"�u>��F�o<�!M��As ȵ�i���E��Q�D�\ҔW�si����Ջ�-���'.F׶��r3椴�բ��;���w��l �<�҂�D(�M��,�]��Z�S#�r��rv��'��3Y\XZ����rR�Z�'��>�fi����~�1"Cy����N�`�m�C*`*gN?g�z����B=�q�r��1V