XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���~�җ �0K�Q+$ѱ2[�na��Oc����-�ގʘ�J[?`��;\>1�H��9Z�A�:��c��o
[���=�酈c����77|�Fhxjmx�2��g�dQ:��)2���jI�����������U"1�8ͅ�.�KN4�@QDO��ġ5�X#Rh�()l[2F����XX3��sO�<_��4�)���؁��/r,�Զ @R�[Ű�k~��WdI��2��>��&a
D+���� �������,r�/g�'���S�=f�%��uǐ���S"
�$]B�:hO,���������X��m��\OaW�E��Tf��9�{6���6ɗ�.��+���#��/�l�J(|�5V+P�*%c)��ZNNf�����x5�h�����"ZT�8�Ik�ܣ-R��$�5pQى;���:1u�k	�)P[�P&&���K�"b�Qܤݯ�.V�@n��k��*���ߑ7`�sv���M�4^=����QF|R���@�$�d�^�����sU��]&PU��U^�zp&��nk�e=�cE���o�~aǝ�j7�23���M
,E'����;N��=Eh}����gε��2���_��x��(�<�ջ8,0���k����N�S� ��Q�g�E˳�a�]�d�����ȥ�\W	K����qxisf[蘒��=���BP<�Om�0l�����Dd�W�)m)���L�˪��$Ǒ>������LVV�����x�>ætűW��.F����M�XlxVHYEB    5e75    1150�?���ұ�zZ��[�g�iS��
�L1��>�o7�S�,�&
�an�Pq��{]kjb�l as��3����,a!>­�t�J��F�J�M���<��eI��W`,������L�}�P����|8�ga�kk�ߑk��v���7.�N�8��b)]����t����b� ��K� ����!T81W���Z�@�"��9_�Q���S`�*���B�T�A����4&o�Pwh�8)�z�Ƴ	\����g �
��w/M�Ls	�V ��A������#���q��p�&mʨ�_o Q"i/���z�;��مL'}�d���� �g�V;�58�b��AT�M�#�w�FFC�F9��w��9r�����:U��S��w�6���?u�#���O�R&�bRt�
;�0@Wl��/����N��^��k�4͌��]tvS��L�����.Ry��Q��a"I�a�)r��Um�w��Ww p%���+#9Suش(��ayw �l"z����k�'��@ ��Ľ6�:��7n5��H�����0�d��T�+�6#R1��)3&�h��(C���/Q�Z�0]��a��~iq	vt�
���vY�X�A�0�}3��6��6L��W�N����������?)})1���7�C����GI'&%N��[�����R���q�ZTPR�5��T�G?�p�q���2�TlupTm=���a�v��T��oל]��!�/���ih�PoA?�]e��G�DTo���t�ƫ����T�*I��T �2��S� 逬�n�ݓ�J�g�َ1</�f[@���䜲u��AL�BT1�"T�\k�������e��l����Ԝ��� �yhyL.��5�����q��m����=r9�U�Ic���է�N��5�sc�$0���-��#��b� Z�*�m[�"Y��7yCOҋ�cKy0};KL�hY����.)6�Q�\�z�І�f ���v�2��z|%��*#����f(�O`�*��=ilN?%�S�2�����:�/��h����7I.9_/���I��'.���h���P+=H��'�� ~B�Xj}*�����@,�fҺ�ݧX�E�-��PNeԥ�S��!������]#7-�1����99�F���0�0Z����	m��&p�g��-\��@�]B��z	 ה���y�-�i8ϛ>2@�Mx�w�m�;�x���H̭�-X#)��-�@
`��{5<xp���	���������(%��i�g�N�Cq0aD�M�%	��	���^��I�tM|���G�J�`VyIҡ�&qa>�m�U"�9��Pe*���-S�V1D�����Z̛)O%����^�>]U�f-0T���,����6���e���S47x�n�y	�|�����ֳ��Vp����.�6?ù%�J���jC����1����0$�K����tܬ�$�w��i`�G�F���I��ȩը�r-��E����-�=:l��c~˄�Y�Q���k�*���a�XJR�~���;�[~������*��I��D$L�@Q9�؃�<���#�x�[m�.�{�������Ko��kw�_=s	��D���7T"ˑf��]3����\-r/�%�q,�ch}>
�&�԰6���7Ee�n̫�j���W�'��"�~o�ch\d�?7�_�{����="�T#��v]���>J��7�Ǟ&�����h^�~*+�q�@��1(fr�ݹ�j�U=dY[�u�H)5��J7Io4Lh璖o"łbm�zf�DS�r�+h7�H��Ya=$
0��U����
�;!�rfR>7�S='����'��+�'h���+�oa�����[d.@s�}G�Q|��D�r�r�_S��s=Y��M���^�&��^��.v�m��a�}{u;�2������s�0+��j����r�)�}j.��X"Ⱦc�Z��^��DEG�At6��'���64t�<���O�%��bdY����5糗$�@��y թ��P���Jr�<U���ã��D]mۏV��f�J�	t�\D,�-kՉ�Us��@׷V��t;G8l#�(T�w(�Z>7d��!:-ZG\��>�QR_;KlN<�?P�v{]�Hȇ)�q	�2�W,�H���(�8U^+����)CɁ1w������s�HEQ>ĸ�IM���J�d����$���'4Ze���5�=g�w��wl�E����@蟇X4�&��:�<N�G�tx��aSJ"���7z����l��;�0�e���g�x�o3 �X����${��")��X8ј�U�  NDB�H���a�5;F;4��y{�]"Dk��y_���-D]D75G����!�������]�(��J�3�x엎
w�L09`fzn�j�lzݴO�!�Od�Zw�D��I�l�硻�g_1��3v|w�G�I�Y^�jՀ�.�q�M�y{G�r��7����c�)"Wf��"b5���5J�{_2M4��,��2����h~���L�L��������8ƻ7��w� �N���k�xe@�����2�ֆ2w�!�t��#�l�'aѳQ��6"Bg����_����������������[�"B@3�5��
H��Z�F3��ksf��N�*���h,e��.8Uu��cݨW�uF�|3�\4@�1ׄz�T��}'vY%����K������ sꏀ��=V}��E>��ʐ������ɼ�{��	�G��ngG�b����t(}�Q�	ɵj���ñ-�:���jE��b��"6M)}�� ѳ�l�:�`G��$K�u�eBxI��sS	�Q���]���{�K���8J�+1��$��3r��<�e:�F�O���3���z�@̽GZՕ�#���e�d�^�8~�9Jf�w�a�e��R���'4�4���W�݋G����x�rHw���
V��u���ޝ�՞�<,b�P������Հ,T,&��s)v��[����@���[	����P�h��
��A�pӈ|O!l�s��P�Xe�!JUǿ�f���H�ܪ%���S�V���(�,�n��.�g���3�T��e����jk�t1��lA��b��O�y�y��X�ݠI����(�� ���7��n�vp��wg��<�QLgt3��m��
��p�?�{�G��B,CKf@Q���8�2z���$�1Վ����Y�;�l��o�X">V��o�\�_��1�/�"�_����Y˂�~��O�
`�Z��.��r��ޮ7��X"ѵ���+xCKr��K^�eh5�C�8�ga�6���I(;1f<k�d�	,��}�M�����[1h�^�E��ڭl����ɿ��� �´�r$��D팖��'�1�X��+�z�)��ꯗt?�%$A�l���zS�
_�R��`�Lkd�J���̔q�ee�[�.ڹ���g�Bd��m>Q�k$s��j��������;�l�p�@���щ���y)�g�E�@WzϷ��R&��+�8S��2��D{������3X�7�㾑�8	 �&¢3I�U���hk����<%Ծ�iZ��������XU~D�Gx�۸?NE�?B�0�&��3y5N5���B�./T�U��0�o�����aߴ4�@!ޗЊ�/A�ч�epB 6�T>��/�r8���	8eI]��	��C��a$��r�T;Z�&�	T����:N@�(��RN��ⲉ�t�wA��d���lӈ�16U0]+�Lœ��g5�1-z-�G�x�0$ϱ��xG�8�d�z�9�u
��xːF,���L�v���%�f%e����&}��c��̵�G曑H��V+{p�=$&�9�1�^x�	\҃*��Z���S!�eej��̰9h'���l�&{㖡���ɅMj-"�}m���GGCخS�f2Xu�N�s����g�`}nA� &9����9���F)SQ��ȍ�a�3���i�{��M�[N��+�Gb!�uPM�\Y�1�z
���*N�n^麍���m��|0hiTO�ߟ\
,KN�r���+�#��!��7���+s�fì����M�<���9W �A(VWǍ�R3M�]ˣ��E\�I��nOǇ�ܐ�C��zd�ֲ�P<zM;K2���ߢ��h{����\�ܷ����ٕ����HD{î����v��0����T��f`�� �֦��-omQU�;��w�I&�m��Tu��\�����!��ž
fI��!@���w~�
��V���菽f;�'�蹍H�^��'c�U�nL��r�)sWلupT�}���AS6�V	�}o7�J�@,O���r ��)�Nv�$u$�z�@�&5�r5��RY�?2�Y�48��_�.T��0ȝو���k���q`=���� �f�Y���x��lz(@�񓺱�iX