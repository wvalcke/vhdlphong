XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����1�V�A"WF��pB�����%��~���/=��yP�����K>t�y�L!�(q�n�UH��)pv\�2��m�-r��!���$=]�\�Պ�c�bc�/C�q_3K���&�9R����%��AmԹ���h�'���Z��f}���Y�m̧V(bl5ZN�.^N�� 6��'���aw�a9�E�A"W��wn��ֳ���,���A������~���R6�l�
�h%��# �s�c�X�|��Q��&��ƺ�݄5�hpR"Y����Bi]��G�g�s����}��k%o B�:�("����7V��_���A'sۡ�$v����݃�褝�ݪ�f�_1ј+0eF[\K2qΈ�z骆>ա�Gߕ�"���D �������m�]�ܨ�D6=����+X[׻8W)c�Jir�ɯ�rYI:p��0�����vO�Jw+Aʏ�$��l���R�
U��e��G>�A�L��@�T�J~e1=�}�dxg��@�S�E]~JR�Z��Q��@e�.�YyL>o�`��hq �aHr:1.�:]�`���p��;t�4�p�]�(r�`IńZ&FK���	,�шn�����Q����V��Pu����M`��W(7t:>!�J� b	q�$Q8���@���SZ�s�E�x?�����G'Q������o�%Ip���,l��i�����'���!z���jO[�����,q��
�QB�rC"�?5.S���k��T<�F�u
�����o8�G#�֛؉�?4wA��gї�*XlxVHYEB    1795     7b0"n^�Z̈́��(�nk��w���#�)�YV�*��Y�:�Qo�o�̝:�f�"r���A!�Q+�2Rr�n2!��+�nT�^`N�Kԝ��Xl��2���[�ϊ]��t�=��W���hK�YA
F��\�?�kL�������i��\��YO��<���C�úI��_��C��-��{E�5Ꮆ���yDKHazGjx4\�B�Zl"U�.6������b�4H�E�-ZJ@t��U�x<�D�)K�@8ךN;��m�.��^"�ܮ��������ku�!�]8�ͺO?�e%s��� g@E�8��T�2�Ě2��9�P�F���������LT6�j�ڹ��3eh	�K����{y.��O`$�L,��NNB�V���
P~�ɱɜ��"�,3��R��e>��|C�{).6���Vbp��<t����i���J���4d�_��=��4� �r����#���ۑ9{c�O��*@���Pb�?5����U�wp�eʫ��;�;��MGX��\g����g��$��Y̓#��X�/����qyV��W�]�n&k�
����:�thT
�44)M� �R@&���`��և�4�����׻G��/�:憶��5��LȨ�5��=���S��bt��k���41�g+C� W�{!�v�d��X���3���	�y�Ծ}C;��]V�c����o��n�k�	\>� �}�g����9ls���kL쏗���?�����|m�k` �����:ٶ+n���KB ��F��N� �K[1�q�U/�����n\��K��)}���c�b�U��3�>'էN$�RE��l��٭-�R�R�C߈ÎcRls�Q�Հ�Qp� }f�k����7���e�<(�h���)$�0���A�6h���3cV�w���g�
{b��B�D���#_ɬ�ɶ6P�S�;=��BT�ZC"w��Sqv�P��.=[�t�8�cT�i�1���һ��tL�j��h���.�{�$�k@�W�m��DW��yc��µ�`��S�Ɲ@������-�j'#؛�6uˈsI���8&��-�aB�pU+.$���t\�������C��uz��=�Z��{1����/���:�L^��5�*m{�������R����= ��q�eV�E^��7��
vEɇ�L$�S A�`� T�N��zx����b}ҫ#�y?D��]>���}����{q�	Es���\b�&:V*��ښ�
���//
z܀�������un�y��\G~̒
6��|m'L��]����rjQ�3�)�߿�	�|�姸r�	-��
��X{��
o��r�⠎yT��_���,i4�ȋ�I�((���@Ћ��e#���zŃ��g�ۜ0���X,;i���G�/�5Fd�.�C��d�e���F�k�0>����S�\./�m!� ��<�n�j��-:�o�T�������v� ��w�$Sc~�2D�	j16.�Tf�A,�4Kk�p�<b&\�H"��zG��o���<~gs{MU��o��[V������%��>�T���ʳ$�S�����@�r�����p �@�`X,J�m��27��L�	���ߙ�$>�
�D�ȄcY �ގ��:\�vX�TÀ����&$~d��+��}�'@+�d�M�Z̹ЮCr����V���0�0[>ye�A����8���inտ�(C}�o�W1H��7IC��mE;����gkp�v��h΢�5f����/�:�B�/���[�/8����y�(Q��>�0|i
�i!�8Tp?��R��+�D%��@0F%\���Ճ�S-��z�,mV��8_�P\S	i#�5%���(煓y�����!�q5��IAB 0�I��$:�]6��\���Ӧħ!�8D�b���������]v�B�J6���*l��`�QidkzX>%ԌWׄ_��<-7:���~&̷�